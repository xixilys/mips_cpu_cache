module alu(
  input  [23:0] io_ctrl,
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_result,
  output        io_overflow
);
  wire [4:0] sa = io_in1[4:0]; // @[alu.scala 22:28]
  wire [31:0] answer_and = io_in1 & io_in2; // @[alu.scala 24:32]
  wire [31:0] answer_or = io_in1 | io_in2; // @[alu.scala 25:32]
  wire [31:0] answer_xor = io_in1 ^ io_in2; // @[alu.scala 26:32]
  wire [31:0] answer_nor = ~answer_or; // @[alu.scala 27:25]
  wire  answer_slt = $signed(io_in1) < $signed(io_in2); // @[alu.scala 29:43]
  wire  answer_sltu = io_in1 < io_in2; // @[alu.scala 30:36]
  wire [62:0] _GEN_5 = {{31'd0}, io_in2}; // @[alu.scala 31:31]
  wire [62:0] answer_sll = _GEN_5 << sa; // @[alu.scala 31:31]
  wire [31:0] answer_srl = io_in2 >> sa; // @[alu.scala 33:31]
  wire [31:0] answer_sra = $signed(io_in2) >>> sa; // @[alu.scala 34:46]
  wire [31:0] answer_lui = {io_in2[15:0],16'h0}; // @[Cat.scala 31:58]
  wire [32:0] in1_extend = {io_in1[31],io_in1}; // @[Cat.scala 31:58]
  wire [32:0] in2_extend = {io_in2[31],io_in2}; // @[Cat.scala 31:58]
  wire [32:0] answer_add = in1_extend + in2_extend; // @[alu.scala 41:35]
  wire [32:0] answer_sub = in1_extend - in2_extend; // @[alu.scala 42:35]
  wire [31:0] _io_result_T_22 = io_ctrl[1] ? answer_add[31:0] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_23 = io_ctrl[2] ? answer_add[31:0] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_24 = io_ctrl[3] ? answer_add[31:0] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_25 = io_ctrl[17] ? answer_sub[31:0] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_26 = io_ctrl[18] ? answer_sub[31:0] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_27 = io_ctrl[19] ? answer_sub[31:0] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_28 = io_ctrl[4] ? answer_and : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_29 = io_ctrl[11] ? answer_or : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_30 = io_ctrl[10] ? answer_nor : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_31 = io_ctrl[20] ? answer_xor : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_32 = io_ctrl[7] ? answer_lui : 32'h0; // @[Mux.scala 27:73]
  wire [62:0] _io_result_T_33 = io_ctrl[12] ? answer_sll : 63'h0; // @[Mux.scala 27:73]
  wire  _io_result_T_34 = io_ctrl[13] & answer_slt; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_35 = io_ctrl[15] ? answer_sra : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_36 = io_ctrl[16] ? answer_srl : 32'h0; // @[Mux.scala 27:73]
  wire  _io_result_T_37 = io_ctrl[14] & answer_sltu; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_38 = _io_result_T_22 | _io_result_T_23; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_39 = _io_result_T_38 | _io_result_T_24; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_40 = _io_result_T_39 | _io_result_T_25; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_41 = _io_result_T_40 | _io_result_T_26; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_42 = _io_result_T_41 | _io_result_T_27; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_43 = _io_result_T_42 | _io_result_T_28; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_44 = _io_result_T_43 | _io_result_T_29; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_45 = _io_result_T_44 | _io_result_T_30; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_46 = _io_result_T_45 | _io_result_T_31; // @[Mux.scala 27:73]
  wire [31:0] _io_result_T_47 = _io_result_T_46 | _io_result_T_32; // @[Mux.scala 27:73]
  wire [62:0] _GEN_0 = {{31'd0}, _io_result_T_47}; // @[Mux.scala 27:73]
  wire [62:0] _io_result_T_48 = _GEN_0 | _io_result_T_33; // @[Mux.scala 27:73]
  wire [62:0] _GEN_1 = {{62'd0}, _io_result_T_34}; // @[Mux.scala 27:73]
  wire [62:0] _io_result_T_49 = _io_result_T_48 | _GEN_1; // @[Mux.scala 27:73]
  wire [62:0] _GEN_2 = {{31'd0}, _io_result_T_35}; // @[Mux.scala 27:73]
  wire [62:0] _io_result_T_50 = _io_result_T_49 | _GEN_2; // @[Mux.scala 27:73]
  wire [62:0] _GEN_3 = {{31'd0}, _io_result_T_36}; // @[Mux.scala 27:73]
  wire [62:0] _io_result_T_51 = _io_result_T_50 | _GEN_3; // @[Mux.scala 27:73]
  wire [62:0] _GEN_4 = {{62'd0}, _io_result_T_37}; // @[Mux.scala 27:73]
  wire [62:0] _io_result_T_52 = _io_result_T_51 | _GEN_4; // @[Mux.scala 27:73]
  assign io_result = _io_result_T_52[31:0]; // @[alu.scala 44:15]
  assign io_overflow = io_ctrl[2] & answer_add[32] != answer_add[31] | io_ctrl[18] & answer_sub[32] != answer_sub[31]; // @[alu.scala 62:79]
endmodule
module br(
  input         reset,
  input  [31:0] io_rs,
  input  [31:0] io_rt,
  input  [5:0]  io_branch,
  output        io_exe
);
  wire  _result_T_1 = $signed(io_rs) < 32'sh0; // @[br.scala 29:38]
  wire  _result_T_3 = $signed(io_rs) <= 32'sh0; // @[br.scala 30:37]
  wire  _result_T_5 = $signed(io_rs) > 32'sh0; // @[br.scala 31:37]
  wire  _result_T_7 = $signed(io_rs) >= 32'sh0; // @[br.scala 32:37]
  wire  _result_T_8 = io_rs != io_rt; // @[br.scala 33:30]
  wire  _result_T_9 = io_rs == io_rt; // @[br.scala 34:30]
  wire [5:0] result = {_result_T_1,_result_T_3,_result_T_5,_result_T_7,_result_T_8,_result_T_9}; // @[Cat.scala 31:58]
  wire [5:0] _io_exe_T_4 = result & io_branch; // @[br.scala 35:57]
  assign io_exe = ~reset & _io_exe_T_4 != 6'h0; // @[br.scala 35:45]
endmodule
module cfu(
  input        reset,
  input        io_Inst_Fifo_Empty,
  input        io_dmem_calD,
  input        io_BranchD_Flag,
  input        io_JRD,
  input        io_CanBranchD,
  input        io_DivPendingE,
  input        io_DataPendingM,
  input        io_InException,
  input  [4:0] io_WriteRegE,
  input        io_RegWriteE,
  input  [1:0] io_HiLoToRegE,
  input        io_CP0ToRegE,
  input  [4:0] io_WriteRegM,
  input        io_MemToRegM,
  input        io_RegWriteM,
  input  [1:0] io_HiLoWriteM,
  input        io_CP0WriteM,
  input  [4:0] io_WriteRegM2,
  input        io_MemToRegM2,
  input        io_RegWriteM2,
  input  [1:0] io_HiLoWriteM2,
  input        io_CP0WriteM2,
  input  [4:0] io_WriteRegW,
  input        io_RegWriteW,
  input  [1:0] io_HiLoWriteW,
  input        io_CP0WriteW,
  input  [4:0] io_ReadCP0AddrE,
  input  [2:0] io_ReadCP0SelE,
  input  [4:0] io_WriteCP0AddrM,
  input  [2:0] io_WriteCP0SelM,
  input  [4:0] io_WriteCP0AddrM2,
  input  [2:0] io_WriteCP0SelM2,
  input  [4:0] io_RsD,
  input  [4:0] io_RtD,
  input  [4:0] io_RsE,
  input  [4:0] io_RtE,
  output       io_StallF,
  output       io_StallD,
  output       io_StallE,
  output       io_StallM,
  output       io_StallM2,
  output       io_StallW,
  output       io_FlushD,
  output       io_FlushE,
  output       io_FlushM,
  output       io_FlushM2,
  output       io_FlushW,
  output [1:0] io_ForwardAE,
  output [1:0] io_ForwardBE,
  output [1:0] io_ForwardAD,
  output [1:0] io_ForwardBD,
  output [1:0] io_ForwardHE,
  output [1:0] io_ForwardCP0E
);
  wire  _io_ForwardAD_T_3 = io_RsD == io_WriteRegM & io_RegWriteM; // @[cfu.scala 107:73]
  wire  _io_ForwardAD_T_5 = ~io_MemToRegM; // @[cfu.scala 107:99]
  wire  _io_ForwardAD_T_9 = io_RsD == io_WriteRegM2 & io_RegWriteM2; // @[cfu.scala 108:34]
  wire  _io_ForwardAD_T_11 = ~io_MemToRegM2; // @[cfu.scala 108:61]
  wire  _io_ForwardAD_T_12 = io_RsD == io_WriteRegM2 & io_RegWriteM2 & ~io_MemToRegM2; // @[cfu.scala 108:58]
  wire [1:0] _io_ForwardAD_T_13 = _io_ForwardAD_T_12 ? 2'h2 : 2'h0; // @[cfu.scala 107:131]
  wire [1:0] _io_ForwardAD_T_14 = io_RsD == io_WriteRegM & io_RegWriteM & ~io_MemToRegM ? 2'h1 : _io_ForwardAD_T_13; // @[cfu.scala 107:48]
  wire  _io_ForwardBD_T_3 = io_RtD == io_WriteRegM & io_RegWriteM; // @[cfu.scala 109:73]
  wire  _io_ForwardBD_T_9 = io_RtD == io_WriteRegM2 & io_RegWriteM2; // @[cfu.scala 110:34]
  wire  _io_ForwardBD_T_12 = io_RtD == io_WriteRegM2 & io_RegWriteM2 & _io_ForwardAD_T_11; // @[cfu.scala 110:58]
  wire [1:0] _io_ForwardBD_T_13 = _io_ForwardBD_T_12 ? 2'h2 : 2'h0; // @[cfu.scala 109:131]
  wire [1:0] _io_ForwardBD_T_14 = io_RtD == io_WriteRegM & io_RegWriteM & _io_ForwardAD_T_5 ? 2'h1 : _io_ForwardBD_T_13; // @[cfu.scala 109:48]
  wire  _io_ForwardAE_T_3 = io_RsE == io_WriteRegM & io_RegWriteM; // @[cfu.scala 116:34]
  wire  _io_ForwardAE_T_6 = io_RsE == io_WriteRegM & io_RegWriteM & _io_ForwardAD_T_5; // @[cfu.scala 116:57]
  wire  _io_ForwardAE_T_9 = io_RsE == io_WriteRegM2 & io_RegWriteM2; // @[cfu.scala 117:35]
  wire  _io_ForwardAE_T_12 = io_RsE == io_WriteRegM2 & io_RegWriteM2 & _io_ForwardAD_T_11; // @[cfu.scala 117:59]
  wire  _io_ForwardAE_T_15 = io_RsE == io_WriteRegW & io_RegWriteW; // @[cfu.scala 118:34]
  wire [1:0] _io_ForwardAE_T_17 = _io_ForwardAE_T_12 ? 2'h3 : {{1'd0}, _io_ForwardAE_T_15}; // @[Mux.scala 101:16]
  wire [1:0] _io_ForwardAE_T_18 = _io_ForwardAE_T_6 ? 2'h2 : _io_ForwardAE_T_17; // @[Mux.scala 101:16]
  wire  _io_ForwardBE_T_3 = io_RtE == io_WriteRegM & io_RegWriteM; // @[cfu.scala 123:34]
  wire  _io_ForwardBE_T_6 = io_RtE == io_WriteRegM & io_RegWriteM & _io_ForwardAD_T_5; // @[cfu.scala 123:57]
  wire  _io_ForwardBE_T_9 = io_RtE == io_WriteRegM2 & io_RegWriteM2; // @[cfu.scala 124:35]
  wire  _io_ForwardBE_T_12 = io_RtE == io_WriteRegM2 & io_RegWriteM2 & _io_ForwardAD_T_11; // @[cfu.scala 124:59]
  wire  _io_ForwardBE_T_15 = io_RtE == io_WriteRegW & io_RegWriteW; // @[cfu.scala 125:34]
  wire [1:0] _io_ForwardBE_T_17 = _io_ForwardBE_T_12 ? 2'h3 : {{1'd0}, _io_ForwardBE_T_15}; // @[Mux.scala 101:16]
  wire [1:0] _io_ForwardBE_T_18 = _io_ForwardBE_T_6 ? 2'h2 : _io_ForwardBE_T_17; // @[Mux.scala 101:16]
  wire [1:0] _io_ForwardHE_T = io_HiLoToRegE & io_HiLoWriteM; // @[cfu.scala 135:25]
  wire  _io_ForwardHE_T_1 = _io_ForwardHE_T != 2'h0; // @[cfu.scala 135:42]
  wire [1:0] _io_ForwardHE_T_2 = io_HiLoToRegE & io_HiLoWriteM2; // @[cfu.scala 136:25]
  wire  _io_ForwardHE_T_3 = _io_ForwardHE_T_2 != 2'h0; // @[cfu.scala 136:43]
  wire [1:0] _io_ForwardHE_T_4 = io_HiLoToRegE & io_HiLoWriteW; // @[cfu.scala 137:25]
  wire  _io_ForwardHE_T_5 = _io_ForwardHE_T_4 != 2'h0; // @[cfu.scala 137:42]
  wire [1:0] _io_ForwardHE_T_7 = _io_ForwardHE_T_3 ? 2'h3 : {{1'd0}, _io_ForwardHE_T_5}; // @[Mux.scala 101:16]
  wire [5:0] _io_ForwardCP0E_T_2 = {io_ReadCP0AddrE,io_ReadCP0SelE[0]}; // @[Cat.scala 31:58]
  wire [5:0] _io_ForwardCP0E_T_4 = {io_WriteCP0AddrM,io_WriteCP0SelM[0]}; // @[Cat.scala 31:58]
  wire  _io_ForwardCP0E_T_7 = _io_ForwardCP0E_T_2 == _io_ForwardCP0E_T_4 & io_CP0WriteM; // @[cfu.scala 141:96]
  wire [5:0] _io_ForwardCP0E_T_11 = {io_WriteCP0AddrM2,io_WriteCP0SelM2[0]}; // @[Cat.scala 31:58]
  wire  _io_ForwardCP0E_T_14 = _io_ForwardCP0E_T_2 == _io_ForwardCP0E_T_11 & io_CP0WriteM2; // @[cfu.scala 142:98]
  wire [1:0] _io_ForwardCP0E_T_15 = _io_ForwardCP0E_T_14 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _io_ForwardCP0E_T_16 = _io_ForwardCP0E_T_7 ? 2'h1 : _io_ForwardCP0E_T_15; // @[Mux.scala 101:16]
  wire  _br_Stall_T_4 = io_WriteRegE == io_RsD; // @[cfu.scala 154:48]
  wire  _br_Stall_T_9 = io_WriteRegM == io_RsD; // @[cfu.scala 155:47]
  wire  _br_Stall_T_12 = io_MemToRegM & (io_WriteRegM == io_RsD | io_WriteRegM == io_RtD); // @[cfu.scala 155:30]
  wire  _br_Stall_T_13 = io_RegWriteE & (io_WriteRegE == io_RsD | io_WriteRegE == io_RtD) | _br_Stall_T_12; // @[cfu.scala 154:88]
  wire  _br_Stall_T_15 = io_WriteRegM2 == io_RsD; // @[cfu.scala 156:49]
  wire  _br_Stall_T_18 = io_MemToRegM2 & (io_WriteRegM2 == io_RsD | io_WriteRegM2 == io_RtD); // @[cfu.scala 156:31]
  wire  _br_Stall_T_19 = _br_Stall_T_13 | _br_Stall_T_18; // @[cfu.scala 155:87]
  wire  _br_Stall_T_20 = io_CanBranchD & io_BranchD_Flag & _br_Stall_T_19; // @[cfu.scala 153:71]
  wire  _br_Stall_T_22 = ~io_InException; // @[cfu.scala 156:95]
  wire  br_Stall = _br_Stall_T_20 & ~io_InException; // @[cfu.scala 156:92]
  wire  _jr_Stall_T_8 = io_MemToRegM & _br_Stall_T_9; // @[cfu.scala 159:30]
  wire  _jr_Stall_T_9 = io_RegWriteE & _br_Stall_T_4 | _jr_Stall_T_8; // @[cfu.scala 158:61]
  wire  _jr_Stall_T_12 = io_MemToRegM2 & _br_Stall_T_15; // @[cfu.scala 160:31]
  wire  _jr_Stall_T_13 = _jr_Stall_T_9 | _jr_Stall_T_12; // @[cfu.scala 159:62]
  wire  _jr_Stall_T_14 = (io_JRD | io_dmem_calD) & _jr_Stall_T_13; // @[cfu.scala 157:60]
  wire  dmem_addr_cal_Stall = _jr_Stall_T_14 & _br_Stall_T_22; // @[cfu.scala 160:65]
  wire  cp0Stall = io_CP0WriteM & io_CP0ToRegE | io_CP0WriteW & io_CP0ToRegE; // @[cfu.scala 168:66]
  wire  _mem2regM_Stall_T_9 = _io_ForwardBE_T_3 & io_MemToRegM; // @[cfu.scala 173:87]
  wire  _mem2regM_Stall_T_10 = _io_ForwardAE_T_3 & io_MemToRegM | _mem2regM_Stall_T_9; // @[cfu.scala 172:120]
  wire  _mem2regM_Stall_T_15 = _io_ForwardAD_T_3 & io_MemToRegM; // @[cfu.scala 174:87]
  wire  _mem2regM_Stall_T_16 = _mem2regM_Stall_T_10 | _mem2regM_Stall_T_15; // @[cfu.scala 173:111]
  wire  _mem2regM_Stall_T_21 = _io_ForwardBD_T_3 & io_MemToRegM; // @[cfu.scala 175:87]
  wire  _mem2regM_Stall_T_22 = _mem2regM_Stall_T_16 | _mem2regM_Stall_T_21; // @[cfu.scala 174:111]
  wire  _mem2regM_Stall_T_27 = _io_ForwardAE_T_9 & io_MemToRegM2; // @[cfu.scala 176:89]
  wire  _mem2regM_Stall_T_28 = _mem2regM_Stall_T_22 | _mem2regM_Stall_T_27; // @[cfu.scala 175:111]
  wire  _mem2regM_Stall_T_33 = _io_ForwardBE_T_9 & io_MemToRegM2; // @[cfu.scala 177:89]
  wire  _mem2regM_Stall_T_34 = _mem2regM_Stall_T_28 | _mem2regM_Stall_T_33; // @[cfu.scala 176:114]
  wire  _mem2regM_Stall_T_39 = _io_ForwardAD_T_9 & io_MemToRegM2; // @[cfu.scala 178:89]
  wire  _mem2regM_Stall_T_40 = _mem2regM_Stall_T_34 | _mem2regM_Stall_T_39; // @[cfu.scala 177:114]
  wire  _mem2regM_Stall_T_45 = _io_ForwardBD_T_9 & io_MemToRegM2; // @[cfu.scala 179:89]
  wire  mem2regM_Stall = _mem2regM_Stall_T_40 | _mem2regM_Stall_T_45; // @[cfu.scala 178:114]
  wire  _has_Stall_T = br_Stall | dmem_addr_cal_Stall; // @[cfu.scala 186:44]
  wire  _io_StallF_T_5 = _has_Stall_T | io_DivPendingE | cp0Stall | io_DataPendingM | mem2regM_Stall; // @[cfu.scala 190:133]
  wire  _io_StallM_T_1 = ~io_DataPendingM; // @[cfu.scala 193:39]
  assign io_StallF = reset | ~(_has_Stall_T | io_DivPendingE | cp0Stall | io_DataPendingM | mem2regM_Stall |
    io_Inst_Fifo_Empty); // @[cfu.scala 190:21]
  assign io_StallD = reset | ~_io_StallF_T_5; // @[cfu.scala 191:21]
  assign io_StallE = reset | ~(io_DivPendingE | cp0Stall | io_DataPendingM | mem2regM_Stall); // @[cfu.scala 192:21]
  assign io_StallM = reset | ~io_DataPendingM; // @[cfu.scala 193:21]
  assign io_StallM2 = reset | _io_StallM_T_1; // @[cfu.scala 194:22]
  assign io_StallW = reset | _io_StallM_T_1; // @[cfu.scala 195:21]
  assign io_FlushD = reset ? 1'h0 : io_InException; // @[cfu.scala 197:21]
  assign io_FlushE = reset ? 1'h0 : io_StallE & _has_Stall_T | io_InException; // @[cfu.scala 198:21]
  assign io_FlushM = reset ? 1'h0 : io_StallM & (cp0Stall | io_DivPendingE | mem2regM_Stall) | io_InException; // @[cfu.scala 199:21]
  assign io_FlushM2 = reset ? 1'h0 : io_InException; // @[cfu.scala 200:22]
  assign io_FlushW = reset ? 1'h0 : io_StallW & (io_DataPendingM | io_InException); // @[cfu.scala 201:21]
  assign io_ForwardAE = io_RsE == 5'h0 ? 2'h0 : _io_ForwardAE_T_18; // @[cfu.scala 115:24]
  assign io_ForwardBE = io_RtE == 5'h0 ? 2'h0 : _io_ForwardBE_T_18; // @[cfu.scala 122:24]
  assign io_ForwardAD = io_RsD == 5'h0 ? 2'h0 : _io_ForwardAD_T_14; // @[cfu.scala 107:24]
  assign io_ForwardBD = io_RtD == 5'h0 ? 2'h0 : _io_ForwardBD_T_14; // @[cfu.scala 109:24]
  assign io_ForwardHE = _io_ForwardHE_T_1 ? 2'h2 : _io_ForwardHE_T_7; // @[Mux.scala 101:16]
  assign io_ForwardCP0E = io_CP0ToRegE ? _io_ForwardCP0E_T_16 : 2'h0; // @[cfu.scala 140:26]
endmodule
module cp0(
  input         clock,
  input         reset,
  input  [4:0]  io_cp0_read_addr,
  input  [2:0]  io_cp0_read_sel,
  input  [4:0]  io_cp0_write_addr,
  input  [2:0]  io_cp0_write_sel,
  input  [31:0] io_cp0_write_data,
  input         io_cp0_write_en,
  input  [5:0]  io_int_i,
  output        io_timer_int_has,
  input  [31:0] io_pc,
  input  [31:0] io_mem_bad_vaddr,
  input  [31:0] io_exception_type_i,
  input         io_in_delayslot,
  input  [1:0]  io_in_branchjump_jr,
  output [31:0] io_return_pc,
  output        io_exception,
  output [31:0] io_cp0_read_data,
  output [31:0] io_epc,
  output [5:0]  io_cp0_status,
  output        io_Int_able,
  output [7:0]  io_asid,
  output [18:0] io_cp0_tlb_read_data_vaddr,
  output [7:0]  io_cp0_tlb_read_data_asid,
  output        io_cp0_tlb_read_data_g,
  output [19:0] io_cp0_tlb_read_data_paddr_0,
  output [19:0] io_cp0_tlb_read_data_paddr_1,
  output [2:0]  io_cp0_tlb_read_data_c_0,
  output [2:0]  io_cp0_tlb_read_data_c_1,
  output        io_cp0_tlb_read_data_d_0,
  output        io_cp0_tlb_read_data_d_1,
  output        io_cp0_tlb_read_data_v_0,
  output        io_cp0_tlb_read_data_v_1,
  input  [18:0] io_cp0_tlb_write_data_vaddr,
  input  [7:0]  io_cp0_tlb_write_data_asid,
  input         io_cp0_tlb_write_data_g,
  input  [19:0] io_cp0_tlb_write_data_paddr_0,
  input  [19:0] io_cp0_tlb_write_data_paddr_1,
  input  [2:0]  io_cp0_tlb_write_data_c_0,
  input  [2:0]  io_cp0_tlb_write_data_c_1,
  input         io_cp0_tlb_write_data_d_0,
  input         io_cp0_tlb_write_data_d_1,
  input         io_cp0_tlb_write_data_v_0,
  input         io_cp0_tlb_write_data_v_1,
  input         io_cp0_tlb_write_en,
  input         io_cp0_index_tlb_write_able
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] cp0_index; // @[cp0.scala 46:28]
  reg [31:0] cp0_random; // @[cp0.scala 47:29]
  reg [31:0] cp0_entrylo0; // @[cp0.scala 48:31]
  reg [31:0] cp0_entrylo1; // @[cp0.scala 49:31]
  reg [31:0] cp0_badvaddr; // @[cp0.scala 51:31]
  reg [31:0] cp0_count; // @[cp0.scala 52:28]
  reg [31:0] cp0_entryhi; // @[cp0.scala 53:30]
  reg [31:0] cp0_compare; // @[cp0.scala 54:30]
  reg [31:0] cp0_status; // @[cp0.scala 55:29]
  reg [31:0] cp0_cause; // @[cp0.scala 56:28]
  reg [31:0] cp0_epc; // @[cp0.scala 57:26]
  reg [31:0] cp0_ebase; // @[cp0.scala 60:28]
  reg [31:0] cp0_config0; // @[cp0.scala 61:30]
  reg  cp0_counter_half; // @[cp0.scala 64:35]
  reg [31:0] plus_380_exception_pc; // @[cp0.scala 73:40]
  wire [31:0] _plus_380_exception_pc_T_3 = {cp0_ebase[31:12],12'h180}; // @[Cat.scala 31:58]
  reg [31:0] plus_200_exception_pc; // @[cp0.scala 75:40]
  wire [31:0] _plus_200_exception_pc_T_3 = {cp0_ebase[31:12],12'h0}; // @[Cat.scala 31:58]
  wire  _io_Int_able_T_1 = ~cp0_status[1]; // @[cp0.scala 82:20]
  wire [7:0] _int_signal_T_2 = cp0_status[15:8] & cp0_cause[15:8]; // @[cp0.scala 86:41]
  wire  int_signal = _int_signal_T_2 != 8'h0 & _io_Int_able_T_1 & cp0_status[0]; // @[cp0.scala 86:89]
  wire [31:0] exception_type = {io_exception_type_i[31:1],int_signal}; // @[Cat.scala 31:58]
  wire  commit_exception = exception_type[30:0] != 31'h0 & _io_Int_able_T_1; // @[cp0.scala 90:58]
  wire  commit_in_delayslot = int_signal | commit_exception ? io_in_delayslot : cp0_cause[31]; // @[cp0.scala 91:34]
  wire [31:0] _commit_eret_T_1 = {{20'd0}, exception_type[31:20]}; // @[cp0.scala 92:65]
  wire  _commit_eret_T_3 = ~_commit_eret_T_1[0]; // @[cp0.scala 92:50]
  wire  commit_eret = exception_type[31] & ~_commit_eret_T_1[0]; // @[cp0.scala 92:47]
  wire  _io_exception_T_1 = commit_exception | commit_eret; // @[cp0.scala 93:43]
  wire [31:0] _commit_next_pc_T_3 = io_pc - 32'h4; // @[cp0.scala 97:11]
  wire [31:0] _commit_next_pc_T_6 = io_pc + 32'h4; // @[cp0.scala 97:61]
  wire [31:0] _commit_next_pc_T_7 = io_in_branchjump_jr != 2'h0 ? io_pc : _commit_next_pc_T_6; // @[cp0.scala 97:21]
  wire [31:0] _commit_epc_T_2 = {{31'd0}, exception_type[31]}; // @[cp0.scala 98:74]
  wire [5:0] read_addr_sel = {io_cp0_read_addr,io_cp0_read_sel[0]}; // @[Cat.scala 31:58]
  wire [5:0] write_addr_sel = {io_cp0_write_addr,io_cp0_write_sel[0]}; // @[Cat.scala 31:58]
  wire  write_and_read_same = write_addr_sel == read_addr_sel & io_cp0_write_en; // @[cp0.scala 130:66]
  wire [17:0] _cp0_read_data_Wire_T_45 = write_and_read_same ? io_cp0_write_data[29:12] : cp0_ebase[29:12]; // @[cp0.scala 152:58]
  wire [31:0] _cp0_read_data_Wire_T_47 = {cp0_ebase[31:30],_cp0_read_data_Wire_T_45,cp0_ebase[11:0]}; // @[Cat.scala 31:58]
  wire [2:0] _cp0_read_data_Wire_T_40 = write_and_read_same ? io_cp0_write_data[2:0] : cp0_config0[2:0]; // @[cp0.scala 150:59]
  wire [31:0] _cp0_read_data_Wire_T_41 = {cp0_config0[31:3],_cp0_read_data_Wire_T_40}; // @[Cat.scala 31:58]
  wire [31:0] _cp0_read_data_Wire_T_36 = write_and_read_same ? io_cp0_write_data : cp0_epc; // @[cp0.scala 148:37]
  wire [1:0] _cp0_read_data_Wire_T_33 = write_and_read_same ? io_cp0_write_data[9:8] : cp0_cause[9:8]; // @[cp0.scala 147:58]
  wire [31:0] _cp0_read_data_Wire_T_35 = {cp0_cause[31:10],_cp0_read_data_Wire_T_33,cp0_cause[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _cp0_read_data_Wire_T_28 = {io_cp0_write_data[31:24],1'h0,io_cp0_write_data[22:8],3'h0,io_cp0_write_data[4
    :0]}; // @[Cat.scala 31:58]
  wire [31:0] _cp0_read_data_Wire_T_29 = write_and_read_same ? _cp0_read_data_Wire_T_28 : cp0_status; // @[cp0.scala 144:37]
  wire [31:0] _cp0_read_data_Wire_T_24 = write_and_read_same ? io_cp0_write_data : cp0_compare; // @[cp0.scala 143:37]
  wire [18:0] _cp0_read_data_Wire_T_19 = write_and_read_same ? io_cp0_write_data[31:13] : cp0_entryhi[31:13]; // @[cp0.scala 141:41]
  wire [7:0] _cp0_read_data_Wire_T_22 = write_and_read_same ? io_cp0_write_data[7:0] : cp0_entryhi[7:0]; // @[cp0.scala 142:37]
  wire [31:0] _cp0_read_data_Wire_T_23 = {_cp0_read_data_Wire_T_19,5'h0,_cp0_read_data_Wire_T_22}; // @[Cat.scala 31:58]
  wire [31:0] _cp0_read_data_Wire_T_16 = write_and_read_same ? io_cp0_write_data : cp0_count; // @[cp0.scala 140:37]
  wire [12:0] _cp0_read_data_Wire_T_14 = write_and_read_same ? {{1'd0}, io_cp0_write_data[24:13]} : 13'h0; // @[cp0.scala 138:50]
  wire [19:0] _cp0_read_data_Wire_T_15 = {7'h0,_cp0_read_data_Wire_T_14}; // @[Cat.scala 31:58]
  wire [25:0] _cp0_read_data_Wire_T_11 = write_and_read_same ? io_cp0_write_data[25:0] : cp0_entrylo1[25:0]; // @[cp0.scala 137:50]
  wire [31:0] _cp0_read_data_Wire_T_12 = {6'h0,_cp0_read_data_Wire_T_11}; // @[Cat.scala 31:58]
  wire [25:0] _cp0_read_data_Wire_T_7 = write_and_read_same ? io_cp0_write_data[25:0] : cp0_entrylo0[25:0]; // @[cp0.scala 136:50]
  wire [31:0] _cp0_read_data_Wire_T_8 = {6'h0,_cp0_read_data_Wire_T_7}; // @[Cat.scala 31:58]
  wire [3:0] _cp0_read_data_Wire_T_3 = write_and_read_same ? io_cp0_write_data[3:0] : cp0_index[3:0]; // @[cp0.scala 134:65]
  wire [31:0] _cp0_read_data_Wire_T_4 = {cp0_index[31],27'h0,_cp0_read_data_Wire_T_3}; // @[Cat.scala 31:58]
  wire [31:0] _cp0_read_data_Wire_T_49 = 6'h0 == read_addr_sel ? _cp0_read_data_Wire_T_4 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _cp0_read_data_Wire_T_51 = 6'h2 == read_addr_sel ? cp0_random : _cp0_read_data_Wire_T_49; // @[Mux.scala 81:58]
  wire [31:0] _cp0_read_data_Wire_T_53 = 6'h4 == read_addr_sel ? _cp0_read_data_Wire_T_8 : _cp0_read_data_Wire_T_51; // @[Mux.scala 81:58]
  wire [31:0] _cp0_read_data_Wire_T_55 = 6'h6 == read_addr_sel ? _cp0_read_data_Wire_T_12 : _cp0_read_data_Wire_T_53; // @[Mux.scala 81:58]
  wire [31:0] _cp0_read_data_Wire_T_57 = 6'ha == read_addr_sel ? {{12'd0}, _cp0_read_data_Wire_T_15} :
    _cp0_read_data_Wire_T_55; // @[Mux.scala 81:58]
  wire [31:0] _cp0_read_data_Wire_T_59 = 6'h10 == read_addr_sel ? cp0_badvaddr : _cp0_read_data_Wire_T_57; // @[Mux.scala 81:58]
  wire [31:0] _cp0_read_data_Wire_T_61 = 6'h12 == read_addr_sel ? _cp0_read_data_Wire_T_16 : _cp0_read_data_Wire_T_59; // @[Mux.scala 81:58]
  wire [31:0] _cp0_read_data_Wire_T_63 = 6'h14 == read_addr_sel ? _cp0_read_data_Wire_T_23 : _cp0_read_data_Wire_T_61; // @[Mux.scala 81:58]
  wire [31:0] _cp0_read_data_Wire_T_65 = 6'h16 == read_addr_sel ? _cp0_read_data_Wire_T_24 : _cp0_read_data_Wire_T_63; // @[Mux.scala 81:58]
  wire [31:0] _cp0_read_data_Wire_T_67 = 6'h18 == read_addr_sel ? _cp0_read_data_Wire_T_29 : _cp0_read_data_Wire_T_65; // @[Mux.scala 81:58]
  wire [31:0] _cp0_read_data_Wire_T_69 = 6'h1a == read_addr_sel ? _cp0_read_data_Wire_T_35 : _cp0_read_data_Wire_T_67; // @[Mux.scala 81:58]
  wire [31:0] _cp0_read_data_Wire_T_71 = 6'h1c == read_addr_sel ? _cp0_read_data_Wire_T_36 : _cp0_read_data_Wire_T_69; // @[Mux.scala 81:58]
  wire [31:0] _cp0_read_data_Wire_T_73 = 6'h1e == read_addr_sel ? 32'h0 : _cp0_read_data_Wire_T_71; // @[Mux.scala 81:58]
  wire [31:0] _cp0_read_data_Wire_T_75 = 6'h20 == read_addr_sel ? _cp0_read_data_Wire_T_41 : _cp0_read_data_Wire_T_73; // @[Mux.scala 81:58]
  wire [31:0] _cp0_read_data_Wire_T_77 = 6'h1 == read_addr_sel ? 32'h1e000000 : _cp0_read_data_Wire_T_75; // @[Mux.scala 81:58]
  wire [31:0] cp0_read_data_Wire = 6'h1f == read_addr_sel ? _cp0_read_data_Wire_T_47 : _cp0_read_data_Wire_T_77; // @[Mux.scala 81:58]
  wire [31:0] _return_pc_Wire_T = {{10'd0}, exception_type[31:10]}; // @[cp0.scala 118:24]
  wire [31:0] _return_pc_Wire_T_2 = {{3'd0}, exception_type[31:3]}; // @[cp0.scala 118:51]
  wire [31:0] _return_pc_Wire_T_5 = {{6'd0}, exception_type[31:6]}; // @[cp0.scala 118:87]
  wire  _return_pc_Wire_T_7 = _return_pc_Wire_T[0] | _return_pc_Wire_T_2[0] | _return_pc_Wire_T_5[0]; // @[cp0.scala 118:70]
  wire  _return_pc_Wire_T_13 = _commit_epc_T_2[0] & _commit_eret_T_3; // @[cp0.scala 119:37]
  wire [31:0] _return_pc_Wire_T_14 = _return_pc_Wire_T_13 ? cp0_epc : plus_380_exception_pc; // @[Mux.scala 101:16]
  wire [31:0] _cause_exccode_Wire_T_2 = {{4'd0}, exception_type[31:4]}; // @[cp0.scala 122:24]
  wire  _cause_exccode_Wire_T_6 = _cause_exccode_Wire_T_2[0] | _commit_eret_T_1[0]; // @[cp0.scala 122:38]
  wire [31:0] _cause_exccode_Wire_T_7 = {{5'd0}, exception_type[31:5]}; // @[cp0.scala 123:23]
  wire [31:0] _cause_exccode_Wire_T_9 = {{8'd0}, exception_type[31:8]}; // @[cp0.scala 123:69]
  wire [31:0] _cause_exccode_Wire_T_11 = {{9'd0}, exception_type[31:9]}; // @[cp0.scala 124:23]
  wire [31:0] _cause_exccode_Wire_T_15 = {{12'd0}, exception_type[31:12]}; // @[cp0.scala 125:23]
  wire [31:0] _cause_exccode_Wire_T_21 = {{2'd0}, exception_type[31:2]}; // @[cp0.scala 126:77]
  wire [31:0] _cause_exccode_Wire_T_23 = {{7'd0}, exception_type[31:7]}; // @[cp0.scala 127:23]
  wire [31:0] _cause_exccode_Wire_T_25 = {{1'd0}, exception_type[31:1]}; // @[cp0.scala 127:78]
  wire [2:0] _cause_exccode_Wire_T_28 = _cause_exccode_Wire_T_6 ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _cause_exccode_Wire_T_29 = _cause_exccode_Wire_T_7[0] ? 3'h5 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _cause_exccode_Wire_T_30 = _cause_exccode_Wire_T_9[0] ? 4'h8 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _cause_exccode_Wire_T_31 = _cause_exccode_Wire_T_11[0] ? 4'h9 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _cause_exccode_Wire_T_32 = _return_pc_Wire_T[0] ? 4'ha : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _cause_exccode_Wire_T_33 = _cause_exccode_Wire_T_15[0] ? 4'hc : 4'h0; // @[Mux.scala 27:73]
  wire [1:0] _cause_exccode_Wire_T_34 = _return_pc_Wire_T_2[0] ? 2'h2 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _cause_exccode_Wire_T_35 = _return_pc_Wire_T_5[0] ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _cause_exccode_Wire_T_36 = _cause_exccode_Wire_T_21[0] ? 2'h2 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _cause_exccode_Wire_T_37 = _cause_exccode_Wire_T_23[0] ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _cause_exccode_Wire_T_40 = _cause_exccode_Wire_T_28 | _cause_exccode_Wire_T_29; // @[Mux.scala 27:73]
  wire [3:0] _GEN_20 = {{1'd0}, _cause_exccode_Wire_T_40}; // @[Mux.scala 27:73]
  wire [3:0] _cause_exccode_Wire_T_41 = _GEN_20 | _cause_exccode_Wire_T_30; // @[Mux.scala 27:73]
  wire [3:0] _cause_exccode_Wire_T_42 = _cause_exccode_Wire_T_41 | _cause_exccode_Wire_T_31; // @[Mux.scala 27:73]
  wire [3:0] _cause_exccode_Wire_T_43 = _cause_exccode_Wire_T_42 | _cause_exccode_Wire_T_32; // @[Mux.scala 27:73]
  wire [3:0] _cause_exccode_Wire_T_44 = _cause_exccode_Wire_T_43 | _cause_exccode_Wire_T_33; // @[Mux.scala 27:73]
  wire [3:0] _GEN_21 = {{2'd0}, _cause_exccode_Wire_T_34}; // @[Mux.scala 27:73]
  wire [3:0] _cause_exccode_Wire_T_45 = _cause_exccode_Wire_T_44 | _GEN_21; // @[Mux.scala 27:73]
  wire [3:0] _GEN_22 = {{2'd0}, _cause_exccode_Wire_T_35}; // @[Mux.scala 27:73]
  wire [3:0] _cause_exccode_Wire_T_46 = _cause_exccode_Wire_T_45 | _GEN_22; // @[Mux.scala 27:73]
  wire [3:0] _GEN_23 = {{2'd0}, _cause_exccode_Wire_T_36}; // @[Mux.scala 27:73]
  wire [3:0] _cause_exccode_Wire_T_47 = _cause_exccode_Wire_T_46 | _GEN_23; // @[Mux.scala 27:73]
  wire [3:0] _GEN_24 = {{2'd0}, _cause_exccode_Wire_T_37}; // @[Mux.scala 27:73]
  wire [3:0] _cause_exccode_Wire_T_48 = _cause_exccode_Wire_T_47 | _GEN_24; // @[Mux.scala 27:73]
  wire [3:0] _GEN_25 = {{3'd0}, _cause_exccode_Wire_T_25[0]}; // @[Mux.scala 27:73]
  wire [3:0] _cause_exccode_Wire_T_49 = _cause_exccode_Wire_T_48 | _GEN_25; // @[Mux.scala 27:73]
  wire  cp0_write_able = io_cp0_write_en & write_addr_sel == 6'h0; // @[cp0.scala 155:49]
  wire  _cp0_index_T_2 = io_cp0_index_tlb_write_able ? io_cp0_write_data[31] : cp0_index[31]; // @[cp0.scala 157:25]
  wire [3:0] _cp0_index_T_5 = cp0_write_able ? io_cp0_write_data[3:0] : cp0_index[3:0]; // @[cp0.scala 157:104]
  wire [27:0] cp0_index_hi = {_cp0_index_T_2,27'h0}; // @[Cat.scala 31:58]
  wire [4:0] _cp0_random_T_2 = cp0_random[4:0] + 5'h1; // @[cp0.scala 158:35]
  wire [31:0] _cp0_entrylo0_T_1 = {6'h0,io_cp0_tlb_write_data_paddr_0,io_cp0_tlb_write_data_c_0,
    io_cp0_tlb_write_data_d_0,io_cp0_tlb_write_data_v_0,io_cp0_tlb_write_data_g}; // @[Cat.scala 31:58]
  wire [25:0] _cp0_entrylo0_T_7 = io_cp0_write_en & write_addr_sel == 6'h4 ? io_cp0_write_data[25:0] : cp0_entrylo0[25:0
    ]; // @[cp0.scala 160:64]
  wire [31:0] _cp0_entrylo1_T_1 = {6'h0,io_cp0_tlb_write_data_paddr_1,io_cp0_tlb_write_data_c_1,
    io_cp0_tlb_write_data_d_1,io_cp0_tlb_write_data_v_1,io_cp0_tlb_write_data_g}; // @[Cat.scala 31:58]
  wire [25:0] _cp0_entrylo1_T_7 = io_cp0_write_en & write_addr_sel == 6'h6 ? io_cp0_write_data[25:0] : cp0_entrylo1[25:0
    ]; // @[cp0.scala 162:64]
  wire [31:0] _cp0_count_T_4 = cp0_count + 32'h1; // @[cp0.scala 165:147]
  wire [31:0] _cp0_entryhi_T = {io_cp0_tlb_write_data_vaddr,5'h0,io_cp0_tlb_write_data_asid}; // @[Cat.scala 31:58]
  wire  _cp0_entryhi_T_3 = io_cp0_write_en & write_addr_sel == 6'h14; // @[cp0.scala 167:56]
  wire [18:0] _cp0_entryhi_T_6 = io_cp0_write_en & write_addr_sel == 6'h14 ? io_cp0_write_data[31:13] : cp0_entryhi[31:
    13]; // @[cp0.scala 167:32]
  wire [7:0] _cp0_entryhi_T_12 = _cp0_entryhi_T_3 ? io_cp0_write_data[7:0] : cp0_entryhi[7:0]; // @[cp0.scala 168:28]
  wire [31:0] _cp0_entryhi_T_13 = {_cp0_entryhi_T_6,5'h0,_cp0_entryhi_T_12}; // @[Cat.scala 31:58]
  wire  _cp0_compare_T_2 = io_cp0_write_en & write_addr_sel == 6'h16; // @[cp0.scala 169:48]
  wire [31:0] _cp0_status_T_4 = {cp0_status[31:2],commit_exception,cp0_status[0]}; // @[Cat.scala 31:58]
  wire  _cp0_status_T_7 = io_cp0_write_en & write_addr_sel == 6'h18; // @[cp0.scala 172:33]
  wire [17:0] _cp0_ebase_T_6 = io_cp0_write_en & write_addr_sel == 6'h1f ? io_cp0_write_data[29:12] : cp0_ebase[29:12]; // @[cp0.scala 174:45]
  wire [19:0] cp0_ebase_hi = {cp0_ebase[31:30],_cp0_ebase_T_6}; // @[Cat.scala 31:58]
  wire  cause_write_en = io_cp0_write_en & write_addr_sel == 6'h1a; // @[cp0.scala 178:48]
  wire  _timer_int_T = cp0_compare != 32'h0; // @[cp0.scala 179:39]
  wire  _timer_int_T_1 = cp0_count == cp0_compare; // @[cp0.scala 179:60]
  wire  _timer_int_T_6 = _cp0_compare_T_2 ? 1'h0 : cp0_cause[30]; // @[cp0.scala 179:109]
  wire  timer_int = cp0_compare != 32'h0 & cp0_count == cp0_compare & ~_cp0_compare_T_2 | _timer_int_T_6; // @[cp0.scala 179:26]
  wire [1:0] _cp0_cause_T_2 = cause_write_en ? io_cp0_write_data[9:8] : cp0_cause[9:8]; // @[cp0.scala 183:82]
  wire [4:0] cause_exccode_Wire = {{1'd0}, _cause_exccode_Wire_T_49}; // @[cp0.scala 105:34 121:24]
  wire [4:0] _cp0_cause_T_5 = cp0_status[1] ? cp0_cause[6:2] : cause_exccode_Wire; // @[cp0.scala 184:38]
  wire [9:0] cp0_cause_lo = {_cp0_cause_T_2,1'h0,_cp0_cause_T_5,2'h0}; // @[Cat.scala 31:58]
  wire [21:0] cp0_cause_hi = {commit_in_delayslot,timer_int,14'h0,io_int_i}; // @[Cat.scala 31:58]
  wire  _cp0_epc_T_3 = io_cp0_write_en & write_addr_sel == 6'h1c; // @[cp0.scala 187:32]
  wire [2:0] _cp0_config0_T_6 = io_cp0_write_en & write_addr_sel == 6'h20 ? io_cp0_write_data[2:0] : cp0_config0[2:0]; // @[cp0.scala 189:45]
  assign io_timer_int_has = _timer_int_T & _timer_int_T_1; // @[cp0.scala 180:44]
  assign io_return_pc = _return_pc_Wire_T_7 ? plus_200_exception_pc : _return_pc_Wire_T_14; // @[Mux.scala 101:16]
  assign io_exception = commit_exception | commit_eret; // @[cp0.scala 93:43]
  assign io_cp0_read_data = reset ? 32'h0 : cp0_read_data_Wire; // @[cp0.scala 103:29]
  assign io_epc = cp0_epc; // @[cp0.scala 81:12]
  assign io_cp0_status = cp0_status[15:10]; // @[cp0.scala 83:33]
  assign io_Int_able = ~cp0_status[1] & cp0_status[0]; // @[cp0.scala 82:36]
  assign io_asid = cp0_entryhi[7:0]; // @[cp0.scala 203:26]
  assign io_cp0_tlb_read_data_vaddr = cp0_entryhi[31:13]; // @[cp0.scala 191:49]
  assign io_cp0_tlb_read_data_asid = cp0_entryhi[7:0]; // @[cp0.scala 192:49]
  assign io_cp0_tlb_read_data_g = cp0_entrylo0[0] & cp0_entrylo1[0]; // @[cp0.scala 193:54]
  assign io_cp0_tlb_read_data_paddr_0 = cp0_entrylo0[25:6]; // @[cp0.scala 194:50]
  assign io_cp0_tlb_read_data_paddr_1 = cp0_entrylo1[25:6]; // @[cp0.scala 195:50]
  assign io_cp0_tlb_read_data_c_0 = cp0_entrylo0[5:3]; // @[cp0.scala 196:50]
  assign io_cp0_tlb_read_data_c_1 = cp0_entrylo1[5:3]; // @[cp0.scala 197:50]
  assign io_cp0_tlb_read_data_d_0 = cp0_entrylo0[2]; // @[cp0.scala 198:50]
  assign io_cp0_tlb_read_data_d_1 = cp0_entrylo1[2]; // @[cp0.scala 199:50]
  assign io_cp0_tlb_read_data_v_0 = cp0_entrylo0[1]; // @[cp0.scala 200:50]
  assign io_cp0_tlb_read_data_v_1 = cp0_entrylo1[1]; // @[cp0.scala 201:50]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Cat.scala 31:58]
      cp0_index <= 32'h0;
    end else begin
      cp0_index <= {cp0_index_hi,_cp0_index_T_5};
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[cp0.scala 47:29]
      cp0_random <= 32'h0; // @[cp0.scala 47:29]
    end else begin
      cp0_random <= {{27'd0}, _cp0_random_T_2}; // @[cp0.scala 158:16]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[cp0.scala 159:24]
      cp0_entrylo0 <= 32'h0;
    end else if (io_cp0_tlb_write_en) begin
      cp0_entrylo0 <= _cp0_entrylo0_T_1;
    end else begin
      cp0_entrylo0 <= {{6'd0}, _cp0_entrylo0_T_7};
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[cp0.scala 161:24]
      cp0_entrylo1 <= 32'h0;
    end else if (io_cp0_tlb_write_en) begin
      cp0_entrylo1 <= _cp0_entrylo1_T_1;
    end else begin
      cp0_entrylo1 <= {{6'd0}, _cp0_entrylo1_T_7};
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[cp0.scala 164:30]
      cp0_badvaddr <= 32'h0; // @[cp0.scala 129:30]
    end else if (commit_exception) begin
      if (_commit_eret_T_1[0] & ~_commit_epc_T_2[0]) begin
        cp0_badvaddr <= io_pc;
      end else begin
        cp0_badvaddr <= io_mem_bad_vaddr;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[cp0.scala 165:30]
      cp0_count <= 32'h0;
    end else if (io_cp0_write_en & write_addr_sel == 6'h12) begin // @[cp0.scala 165:117]
      cp0_count <= io_cp0_write_data;
    end else if (cp0_counter_half) begin
      cp0_count <= _cp0_count_T_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[cp0.scala 166:23]
      cp0_entryhi <= 32'h0;
    end else if (io_cp0_tlb_write_en) begin
      cp0_entryhi <= _cp0_entryhi_T;
    end else begin
      cp0_entryhi <= _cp0_entryhi_T_13;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[cp0.scala 169:24]
      cp0_compare <= 32'h0;
    end else if (io_cp0_write_en & write_addr_sel == 6'h16) begin
      cp0_compare <= io_cp0_write_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Mux.scala 101:16]
      cp0_status <= 32'h400000;
    end else if (_io_exception_T_1) begin // @[Mux.scala 101:16]
      cp0_status <= _cp0_status_T_4;
    end else if (_cp0_status_T_7) begin
      cp0_status <= _cp0_read_data_Wire_T_28;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Cat.scala 31:58]
      cp0_cause <= 32'h0;
    end else begin
      cp0_cause <= {cp0_cause_hi,cp0_cause_lo};
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Mux.scala 101:16]
      cp0_epc <= 32'h0; // @[cp0.scala 98:28 96:{31,53} 97:71]
    end else if (commit_exception) begin // @[Mux.scala 101:16]
      if (!(_commit_eret_T_1[0] & _commit_epc_T_2[0])) begin
        if (int_signal) begin
          if (io_in_delayslot) begin
            cp0_epc <= _commit_next_pc_T_3;
          end else begin
            cp0_epc <= _commit_next_pc_T_7;
          end
        end else if (io_in_delayslot) begin
          cp0_epc <= _commit_next_pc_T_3;
        end else begin
          cp0_epc <= io_pc;
        end
      end
    end else if (_cp0_epc_T_3) begin
      cp0_epc <= io_cp0_write_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Cat.scala 31:58]
      cp0_ebase <= 32'haff00000;
    end else begin
      cp0_ebase <= {cp0_ebase_hi,cp0_ebase[11:0]};
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Cat.scala 31:58]
      cp0_config0 <= 32'h80000082;
    end else begin
      cp0_config0 <= {cp0_config0[31:3],_cp0_config0_T_6};
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[cp0.scala 66:28]
      cp0_counter_half <= 1'h0;
    end else if (clock) begin
      cp0_counter_half <= ~cp0_counter_half;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[cp0.scala 74:33]
      plus_380_exception_pc <= 32'hbfc00380;
    end else if (cp0_status[22]) begin
      plus_380_exception_pc <= 32'hbfc00380;
    end else begin
      plus_380_exception_pc <= _plus_380_exception_pc_T_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[cp0.scala 76:33]
      plus_200_exception_pc <= 32'hbfc00200;
    end else if (cp0_status[22]) begin
      plus_200_exception_pc <= 32'hbfc00200;
    end else begin
      plus_200_exception_pc <= _plus_200_exception_pc_T_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cp0_index = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cp0_random = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  cp0_entrylo0 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  cp0_entrylo1 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  cp0_badvaddr = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  cp0_count = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  cp0_entryhi = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  cp0_compare = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  cp0_status = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  cp0_cause = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  cp0_epc = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  cp0_ebase = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  cp0_config0 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  cp0_counter_half = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  plus_380_exception_pc = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  plus_200_exception_pc = _RAND_15[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    cp0_index = 32'h0;
  end
  if (reset) begin
    cp0_random = 32'h0;
  end
  if (reset) begin
    cp0_entrylo0 = 32'h0;
  end
  if (reset) begin
    cp0_entrylo1 = 32'h0;
  end
  if (reset) begin
    cp0_badvaddr = 32'h0;
  end
  if (reset) begin
    cp0_count = 32'h0;
  end
  if (reset) begin
    cp0_entryhi = 32'h0;
  end
  if (reset) begin
    cp0_compare = 32'h0;
  end
  if (reset) begin
    cp0_status = 32'h400000;
  end
  if (reset) begin
    cp0_cause = 32'h0;
  end
  if (reset) begin
    cp0_epc = 32'h0;
  end
  if (reset) begin
    cp0_ebase = 32'haff00000;
  end
  if (reset) begin
    cp0_config0 = 32'h80000082;
  end
  if (reset) begin
    cp0_counter_half = 1'h0;
  end
  if (reset) begin
    plus_380_exception_pc = 32'hbfc00380;
  end
  if (reset) begin
    plus_200_exception_pc = 32'hbfc00200;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cu(
  input         reset,
  input  [31:0] io1_InstrD,
  output        io1_BadInstrD,
  output        io1_BreakD,
  output        io1_SysCallD,
  output        io1_EretD,
  output [2:0]  io1_Tlb_Control,
  output        io1_commit_cache_ins,
  output        io1_dmem_addr_cal,
  output        io_RegWriteD,
  output        io_MemToRegD,
  output        io_MemWriteD,
  output [23:0] io_ALUCtrlD,
  output [1:0]  io_ALUSrcD,
  output [1:0]  io_RegDstD,
  output        io_ImmUnsigned,
  output        io_LinkD,
  output [1:0]  io_HiLoWriteD,
  output [1:0]  io_HiLoToRegD,
  output        io_CP0WriteD,
  output        io_CP0ToRegD,
  output        io_LoadUnsignedD,
  output [1:0]  io_MemWidthD,
  output [1:0]  io_MemRLD
);
  wire [5:0] OpD = io1_InstrD[31:26]; // @[cu.scala 50:25]
  wire [5:0] FunctD = io1_InstrD[5:0]; // @[cu.scala 51:28]
  wire [4:0] RtD = io1_InstrD[20:16]; // @[cu.scala 53:28]
  wire  coD = io1_InstrD[25]; // @[cu.scala 56:25]
  wire [3:0] coD_res = io1_InstrD[24:21]; // @[cu.scala 57:29]
  wire  _io_LinkD_T_9 = 6'h1 == OpD ? 5'h10 == RtD | 5'h11 == RtD : 6'h3 == OpD; // @[Mux.scala 81:58]
  wire [2:0] _ins_id_T_1 = 6'h22 == FunctD ? 3'h5 : 3'h0; // @[Mux.scala 81:58]
  wire [3:0] _ins_id_T_3 = 6'h24 == FunctD ? 4'hf : {{1'd0}, _ins_id_T_1}; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_5 = 6'h25 == FunctD ? 5'h13 : {{1'd0}, _ins_id_T_3}; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_7 = 6'h2a == FunctD ? 5'h7 : _ins_id_T_5; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_9 = 6'h0 == FunctD ? 5'h17 : _ins_id_T_7; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_11 = 6'h2b == FunctD ? 5'h9 : _ins_id_T_9; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_13 = 6'h26 == FunctD ? 5'h15 : _ins_id_T_11; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_15 = 6'h20 == FunctD ? 5'h1 : _ins_id_T_13; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_17 = 6'h21 == FunctD ? 5'h3 : _ins_id_T_15; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_19 = 6'h23 == FunctD ? 5'h6 : _ins_id_T_17; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_21 = 6'h1a == FunctD ? 5'hb : _ins_id_T_19; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_23 = 6'h1b == FunctD ? 5'hc : _ins_id_T_21; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_25 = 6'h18 == FunctD ? 5'hd : _ins_id_T_23; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_27 = 6'h19 == FunctD ? 5'he : _ins_id_T_25; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_29 = 6'h27 == FunctD ? 5'h12 : _ins_id_T_27; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_31 = 6'h4 == FunctD ? 5'h18 : _ins_id_T_29; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_33 = 6'h3 == FunctD ? 5'h19 : _ins_id_T_31; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_35 = 6'h7 == FunctD ? 5'h1a : _ins_id_T_33; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_37 = 6'h2 == FunctD ? 5'h1b : _ins_id_T_35; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_39 = 6'h6 == FunctD ? 5'h1c : _ins_id_T_37; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_41 = 6'h8 == FunctD ? 6'h27 : {{1'd0}, _ins_id_T_39}; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_43 = 6'h9 == FunctD ? 6'h28 : _ins_id_T_41; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_45 = 6'h10 == FunctD ? 6'h29 : _ins_id_T_43; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_47 = 6'h12 == FunctD ? 6'h2a : _ins_id_T_45; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_49 = 6'h11 == FunctD ? 6'h2b : _ins_id_T_47; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_51 = 6'h13 == FunctD ? 6'h2c : _ins_id_T_49; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_53 = 6'hd == FunctD ? 6'h2d : _ins_id_T_51; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_55 = 6'hc == FunctD ? 6'h2e : _ins_id_T_53; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_57 = 6'h34 == FunctD ? 7'h46 : {{1'd0}, _ins_id_T_55}; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_59 = 6'h36 == FunctD ? 7'h48 : _ins_id_T_57; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_61 = 6'h31 == FunctD ? 7'h4c : _ins_id_T_59; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_63 = 6'h30 == FunctD ? 7'h4a : _ins_id_T_61; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_65 = 6'h32 == FunctD ? 7'h4e : _ins_id_T_63; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_67 = 6'h33 == FunctD ? 7'h50 : _ins_id_T_65; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_69 = 6'hf == FunctD ? 7'h52 : _ins_id_T_67; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_71 = 5'hc == RtD ? 7'h47 : 7'h0; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_73 = 5'he == RtD ? 7'h49 : _ins_id_T_71; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_75 = 5'h8 == RtD ? 7'h4b : _ins_id_T_73; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_77 = 5'h9 == RtD ? 7'h4d : _ins_id_T_75; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_79 = 5'ha == RtD ? 7'h4f : _ins_id_T_77; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_81 = 5'hb == RtD ? 7'h51 : _ins_id_T_79; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_83 = 5'h1 == RtD ? 7'h1f : _ins_id_T_81; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_85 = 5'h11 == RtD ? 7'h20 : _ins_id_T_83; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_87 = 5'h0 == RtD ? 7'h23 : _ins_id_T_85; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_89 = 5'h10 == RtD ? 7'h24 : _ins_id_T_87; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_91 = 6'h8 == FunctD ? 7'h40 : 7'h1; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_93 = 6'h1 == FunctD ? 7'h41 : _ins_id_T_91; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_95 = 6'h2 == FunctD ? 7'h42 : _ins_id_T_93; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_97 = 6'h6 == FunctD ? 7'h43 : _ins_id_T_95; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_99 = 6'h18 == FunctD ? 7'h37 : _ins_id_T_97; // @[Mux.scala 81:58]
  wire [4:0] _GEN_0 = {{1'd0}, coD_res}; // @[Mux.scala 81:61]
  wire [5:0] _ins_id_T_101 = 5'h0 == _GEN_0 ? 6'h38 : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_103 = 5'h4 == _GEN_0 ? 6'h39 : _ins_id_T_101; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_105 = ~coD ? {{1'd0}, _ins_id_T_103} : _ins_id_T_99; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_107 = 6'h2 == FunctD ? 6'h3f : 6'h0; // @[Mux.scala 81:58]
  wire [1:0] _ins_id_T_109 = 6'h8 == OpD ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_111 = 6'hc == OpD ? 5'h10 : {{3'd0}, _ins_id_T_109}; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_113 = 6'h9 == OpD ? 5'h4 : _ins_id_T_111; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_115 = 6'ha == OpD ? 5'h8 : _ins_id_T_113; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_117 = 6'hb == OpD ? 5'ha : _ins_id_T_115; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_119 = 6'hf == OpD ? 5'h11 : _ins_id_T_117; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_121 = 6'hd == OpD ? 5'h14 : _ins_id_T_119; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_123 = 6'he == OpD ? 5'h16 : _ins_id_T_121; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_125 = 6'h4 == OpD ? 5'h1d : _ins_id_T_123; // @[Mux.scala 81:58]
  wire [4:0] _ins_id_T_127 = 6'h5 == OpD ? 5'h1e : _ins_id_T_125; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_129 = 6'h7 == OpD ? 6'h21 : {{1'd0}, _ins_id_T_127}; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_131 = 6'h6 == OpD ? 6'h22 : _ins_id_T_129; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_133 = 6'h2 == OpD ? 6'h25 : _ins_id_T_131; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_135 = 6'h3 == OpD ? 6'h26 : _ins_id_T_133; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_137 = 6'h20 == OpD ? 6'h2f : _ins_id_T_135; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_139 = 6'h24 == OpD ? 6'h30 : _ins_id_T_137; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_141 = 6'h21 == OpD ? 6'h31 : _ins_id_T_139; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_143 = 6'h25 == OpD ? 6'h32 : _ins_id_T_141; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_145 = 6'h23 == OpD ? 6'h33 : _ins_id_T_143; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_147 = 6'h28 == OpD ? 6'h34 : _ins_id_T_145; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_149 = 6'h29 == OpD ? 6'h35 : _ins_id_T_147; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_151 = 6'h2b == OpD ? 6'h36 : _ins_id_T_149; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_153 = 6'h22 == OpD ? 6'h3b : _ins_id_T_151; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_155 = 6'h26 == OpD ? 6'h3c : _ins_id_T_153; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_157 = 6'h2a == OpD ? 6'h3d : _ins_id_T_155; // @[Mux.scala 81:58]
  wire [5:0] _ins_id_T_159 = 6'h2e == OpD ? 6'h3e : _ins_id_T_157; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_161 = 6'h2f == OpD ? 7'h44 : {{1'd0}, _ins_id_T_159}; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_163 = 6'h0 == OpD ? _ins_id_T_69 : _ins_id_T_161; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_165 = 6'h1 == OpD ? _ins_id_T_89 : _ins_id_T_163; // @[Mux.scala 81:58]
  wire [6:0] _ins_id_T_167 = 6'h10 == OpD ? _ins_id_T_105 : _ins_id_T_165; // @[Mux.scala 81:58]
  wire [6:0] ins_id = 6'h1c == OpD ? {{1'd0}, _ins_id_T_107} : _ins_id_T_167; // @[Mux.scala 81:58]
  wire  _io1_Tlb_Control_T = ins_id == 7'h40; // @[cu.scala 245:35]
  wire  _io1_Tlb_Control_T_1 = ins_id == 7'h41; // @[cu.scala 245:57]
  wire  _io1_Tlb_Control_T_2 = ins_id == 7'h42; // @[cu.scala 245:80]
  wire [1:0] io1_Tlb_Control_hi = {_io1_Tlb_Control_T,_io1_Tlb_Control_T_1}; // @[Cat.scala 31:58]
  wire [28:0] _get_controls_T_3 = 7'h2 == ins_id ? 29'h2200000 : 29'h0; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_5 = 7'h5 == ins_id ? 29'h2800000 : _get_controls_T_3; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_7 = 7'hf == ins_id ? 29'h2800000 : _get_controls_T_5; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_9 = 7'h13 == ins_id ? 29'h2800000 : _get_controls_T_7; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_11 = 7'h15 == ins_id ? 29'h2800000 : _get_controls_T_9; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_13 = 7'h7 == ins_id ? 29'h2800000 : _get_controls_T_11; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_15 = 7'h17 == ins_id ? 29'h2c00000 : _get_controls_T_13; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_17 = 7'h10 == ins_id ? 29'h2300000 : _get_controls_T_15; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_19 = 7'h1 == ins_id ? 29'h2800000 : _get_controls_T_17; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_21 = 7'h3 == ins_id ? 29'h2800000 : _get_controls_T_19; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_23 = 7'h4 == ins_id ? 29'h2200000 : _get_controls_T_21; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_25 = 7'h6 == ins_id ? 29'h2800000 : _get_controls_T_23; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_27 = 7'h8 == ins_id ? 29'h2200000 : _get_controls_T_25; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_29 = 7'h9 == ins_id ? 29'h2800000 : _get_controls_T_27; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_31 = 7'ha == ins_id ? 29'h2200000 : _get_controls_T_29; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_33 = 7'hb == ins_id ? 29'h600 : _get_controls_T_31; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_35 = 7'hc == ins_id ? 29'h600 : _get_controls_T_33; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_37 = 7'hd == ins_id ? 29'h600 : _get_controls_T_35; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_39 = 7'he == ins_id ? 29'h600 : _get_controls_T_37; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_41 = 7'h11 == ins_id ? 29'h2200000 : _get_controls_T_39; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_43 = 7'h12 == ins_id ? 29'h2800000 : _get_controls_T_41; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_45 = 7'h14 == ins_id ? 29'h2300000 : _get_controls_T_43; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_47 = 7'h16 == ins_id ? 29'h2300000 : _get_controls_T_45; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_49 = 7'h18 == ins_id ? 29'h2800000 : _get_controls_T_47; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_51 = 7'h19 == ins_id ? 29'h2c00000 : _get_controls_T_49; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_53 = 7'h1a == ins_id ? 29'h2800000 : _get_controls_T_51; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_55 = 7'h1b == ins_id ? 29'h2c00000 : _get_controls_T_53; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_57 = 7'h1c == ins_id ? 29'h2800000 : _get_controls_T_55; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_59 = 7'h1d == ins_id ? 29'h4004000 : _get_controls_T_57; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_61 = 7'h1e == ins_id ? 29'h4008000 : _get_controls_T_59; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_63 = 7'h1f == ins_id ? 29'h4010000 : _get_controls_T_61; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_65 = 7'h20 == ins_id ? 29'h7010800 : _get_controls_T_63; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_67 = 7'h21 == ins_id ? 29'h4020000 : _get_controls_T_65; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_69 = 7'h22 == ins_id ? 29'h4040000 : _get_controls_T_67; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_71 = 7'h23 == ins_id ? 29'h4080000 : _get_controls_T_69; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_73 = 7'h24 == ins_id ? 29'h7080800 : _get_controls_T_71; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_75 = 7'h25 == ins_id ? 29'h2000 : _get_controls_T_73; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_77 = 7'h26 == ins_id ? 29'h3002800 : _get_controls_T_75; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_79 = 7'h27 == ins_id ? 29'h3000 : _get_controls_T_77; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_81 = 7'h28 == ins_id ? 29'h2803800 : _get_controls_T_79; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_83 = 7'h29 == ins_id ? 29'h2800100 : _get_controls_T_81; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_85 = 7'h2a == ins_id ? 29'h2800080 : _get_controls_T_83; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_87 = 7'h2b == ins_id ? 29'h400 : _get_controls_T_85; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_89 = 7'h2c == ins_id ? 29'h200 : _get_controls_T_87; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_91 = 7'h2d == ins_id ? 29'h0 : _get_controls_T_89; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_93 = 7'h2e == ins_id ? 29'h0 : _get_controls_T_91; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_95 = 7'h2f == ins_id ? 29'h2200008 : _get_controls_T_93; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_97 = 7'h30 == ins_id ? 29'h220000c : _get_controls_T_95; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_99 = 7'h31 == ins_id ? 29'h2200009 : _get_controls_T_97; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_101 = 7'h32 == ins_id ? 29'h220000d : _get_controls_T_99; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_103 = 7'h33 == ins_id ? 29'h220000a : _get_controls_T_101; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_105 = 7'h34 == ins_id ? 29'h200010 : _get_controls_T_103; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_107 = 7'h35 == ins_id ? 29'h200011 : _get_controls_T_105; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_109 = 7'h36 == ins_id ? 29'h200012 : _get_controls_T_107; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_111 = 7'h37 == ins_id ? 29'h0 : _get_controls_T_109; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_113 = 7'h38 == ins_id ? 29'h2000020 : _get_controls_T_111; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_115 = 7'h39 == ins_id ? 29'h40 : _get_controls_T_113; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_117 = 7'h3d == ins_id ? 29'h10200012 : _get_controls_T_115; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_119 = 7'h3e == ins_id ? 29'h8200012 : _get_controls_T_117; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_121 = 7'h3b == ins_id ? 29'h1220000a : _get_controls_T_119; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_123 = 7'h3c == ins_id ? 29'ha20000a : _get_controls_T_121; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_125 = 7'h3f == ins_id ? 29'h2800000 : _get_controls_T_123; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_127 = 7'h40 == ins_id ? 29'h20 : _get_controls_T_125; // @[Mux.scala 81:58]
  wire [28:0] _get_controls_T_129 = 7'h41 == ins_id ? 29'h20 : _get_controls_T_127; // @[Mux.scala 81:58]
  wire [28:0] get_controls = 7'h42 == ins_id ? 29'h20 : _get_controls_T_129; // @[Mux.scala 81:58]
  wire [2:0] _get_alu_op_T_66 = 7'h1 == ins_id ? 3'h4 : {{2'd0}, 7'h0 == ins_id}; // @[Mux.scala 81:58]
  wire [2:0] _get_alu_op_T_68 = 7'h2 == ins_id ? 3'h4 : _get_alu_op_T_66; // @[Mux.scala 81:58]
  wire [3:0] _get_alu_op_T_70 = 7'h3 == ins_id ? 4'h8 : {{1'd0}, _get_alu_op_T_68}; // @[Mux.scala 81:58]
  wire [3:0] _get_alu_op_T_72 = 7'h4 == ins_id ? 4'h8 : _get_alu_op_T_70; // @[Mux.scala 81:58]
  wire [18:0] _get_alu_op_T_74 = 7'h5 == ins_id ? 19'h40000 : {{15'd0}, _get_alu_op_T_72}; // @[Mux.scala 81:58]
  wire [19:0] _get_alu_op_T_76 = 7'h6 == ins_id ? 20'h80000 : {{1'd0}, _get_alu_op_T_74}; // @[Mux.scala 81:58]
  wire [19:0] _get_alu_op_T_78 = 7'h7 == ins_id ? 20'h2000 : _get_alu_op_T_76; // @[Mux.scala 81:58]
  wire [19:0] _get_alu_op_T_80 = 7'h8 == ins_id ? 20'h2000 : _get_alu_op_T_78; // @[Mux.scala 81:58]
  wire [19:0] _get_alu_op_T_82 = 7'h9 == ins_id ? 20'h4000 : _get_alu_op_T_80; // @[Mux.scala 81:58]
  wire [19:0] _get_alu_op_T_84 = 7'ha == ins_id ? 20'h4000 : _get_alu_op_T_82; // @[Mux.scala 81:58]
  wire [19:0] _get_alu_op_T_86 = 7'hb == ins_id ? 20'h20 : _get_alu_op_T_84; // @[Mux.scala 81:58]
  wire [19:0] _get_alu_op_T_88 = 7'hc == ins_id ? 20'h40 : _get_alu_op_T_86; // @[Mux.scala 81:58]
  wire [19:0] _get_alu_op_T_90 = 7'hd == ins_id ? 20'h100 : _get_alu_op_T_88; // @[Mux.scala 81:58]
  wire [19:0] _get_alu_op_T_92 = 7'he == ins_id ? 20'h200 : _get_alu_op_T_90; // @[Mux.scala 81:58]
  wire [19:0] _get_alu_op_T_94 = 7'hf == ins_id ? 20'h10 : _get_alu_op_T_92; // @[Mux.scala 81:58]
  wire [19:0] _get_alu_op_T_96 = 7'h10 == ins_id ? 20'h10 : _get_alu_op_T_94; // @[Mux.scala 81:58]
  wire [19:0] _get_alu_op_T_98 = 7'h11 == ins_id ? 20'h80 : _get_alu_op_T_96; // @[Mux.scala 81:58]
  wire [19:0] _get_alu_op_T_100 = 7'h12 == ins_id ? 20'h400 : _get_alu_op_T_98; // @[Mux.scala 81:58]
  wire [19:0] _get_alu_op_T_102 = 7'h13 == ins_id ? 20'h800 : _get_alu_op_T_100; // @[Mux.scala 81:58]
  wire [19:0] _get_alu_op_T_104 = 7'h14 == ins_id ? 20'h800 : _get_alu_op_T_102; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_106 = 7'h15 == ins_id ? 21'h100000 : {{1'd0}, _get_alu_op_T_104}; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_108 = 7'h16 == ins_id ? 21'h100000 : _get_alu_op_T_106; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_110 = 7'h17 == ins_id ? 21'h1000 : _get_alu_op_T_108; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_112 = 7'h18 == ins_id ? 21'h1000 : _get_alu_op_T_110; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_114 = 7'h19 == ins_id ? 21'h8000 : _get_alu_op_T_112; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_116 = 7'h1a == ins_id ? 21'h8000 : _get_alu_op_T_114; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_118 = 7'h1b == ins_id ? 21'h10000 : _get_alu_op_T_116; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_120 = 7'h1c == ins_id ? 21'h10000 : _get_alu_op_T_118; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_122 = 7'h1d == ins_id ? 21'h20000 : _get_alu_op_T_120; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_124 = 7'h1e == ins_id ? 21'h20000 : _get_alu_op_T_122; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_126 = 7'h1f == ins_id ? 21'h20000 : _get_alu_op_T_124; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_128 = 7'h20 == ins_id ? 21'h20000 : _get_alu_op_T_126; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_130 = 7'h21 == ins_id ? 21'h20000 : _get_alu_op_T_128; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_132 = 7'h22 == ins_id ? 21'h20000 : _get_alu_op_T_130; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_134 = 7'h23 == ins_id ? 21'h20000 : _get_alu_op_T_132; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_136 = 7'h24 == ins_id ? 21'h20000 : _get_alu_op_T_134; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_138 = 7'h25 == ins_id ? 21'h1 : _get_alu_op_T_136; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_140 = 7'h26 == ins_id ? 21'h1 : _get_alu_op_T_138; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_142 = 7'h27 == ins_id ? 21'h1 : _get_alu_op_T_140; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_144 = 7'h28 == ins_id ? 21'h1 : _get_alu_op_T_142; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_146 = 7'h29 == ins_id ? 21'h1 : _get_alu_op_T_144; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_148 = 7'h2a == ins_id ? 21'h1 : _get_alu_op_T_146; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_150 = 7'h2b == ins_id ? 21'h1 : _get_alu_op_T_148; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_152 = 7'h2c == ins_id ? 21'h1 : _get_alu_op_T_150; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_154 = 7'h2d == ins_id ? 21'h1 : _get_alu_op_T_152; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_156 = 7'h2e == ins_id ? 21'h1 : _get_alu_op_T_154; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_158 = 7'h2f == ins_id ? 21'h2 : _get_alu_op_T_156; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_160 = 7'h30 == ins_id ? 21'h2 : _get_alu_op_T_158; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_162 = 7'h31 == ins_id ? 21'h2 : _get_alu_op_T_160; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_164 = 7'h32 == ins_id ? 21'h2 : _get_alu_op_T_162; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_166 = 7'h33 == ins_id ? 21'h2 : _get_alu_op_T_164; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_168 = 7'h34 == ins_id ? 21'h2 : _get_alu_op_T_166; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_170 = 7'h35 == ins_id ? 21'h2 : _get_alu_op_T_168; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_172 = 7'h36 == ins_id ? 21'h2 : _get_alu_op_T_170; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_174 = 7'h3d == ins_id ? 21'h2 : _get_alu_op_T_172; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_176 = 7'h3e == ins_id ? 21'h2 : _get_alu_op_T_174; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_178 = 7'h3b == ins_id ? 21'h2 : _get_alu_op_T_176; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_180 = 7'h3c == ins_id ? 21'h2 : _get_alu_op_T_178; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_182 = 7'h37 == ins_id ? 21'h1 : _get_alu_op_T_180; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_184 = 7'h38 == ins_id ? 21'h1 : _get_alu_op_T_182; // @[Mux.scala 81:58]
  wire [20:0] _get_alu_op_T_186 = 7'h39 == ins_id ? 21'h1 : _get_alu_op_T_184; // @[Mux.scala 81:58]
  wire [21:0] _get_alu_op_T_188 = 7'h3f == ins_id ? 22'h200000 : {{1'd0}, _get_alu_op_T_186}; // @[Mux.scala 81:58]
  wire [23:0] get_alu_op = {{2'd0}, _get_alu_op_T_188}; // @[cu.scala 337:26 340:16]
  assign io1_BadInstrD = ins_id == 7'h0; // @[cu.scala 241:29]
  assign io1_BreakD = ins_id == 7'h2d; // @[cu.scala 242:29]
  assign io1_SysCallD = ins_id == 7'h2e; // @[cu.scala 243:29]
  assign io1_EretD = ins_id == 7'h37; // @[cu.scala 244:29]
  assign io1_Tlb_Control = {io1_Tlb_Control_hi,_io1_Tlb_Control_T_2}; // @[Cat.scala 31:58]
  assign io1_commit_cache_ins = io1_InstrD == 32'h3fd0021; // @[cu.scala 246:40]
  assign io1_dmem_addr_cal = 6'h2e == OpD | (6'h2a == OpD | (6'h26 == OpD | (6'h22 == OpD | (6'h2b == OpD | (6'h29 ==
    OpD | (6'h28 == OpD | (6'h23 == OpD | (6'h25 == OpD | (6'h21 == OpD | (6'h24 == OpD | 6'h20 == OpD)))))))))); // @[Mux.scala 81:58]
  assign io_RegWriteD = get_controls[25]; // @[cu.scala 251:33]
  assign io_MemToRegD = get_controls[3]; // @[cu.scala 264:34]
  assign io_MemWriteD = get_controls[4]; // @[cu.scala 263:34]
  assign io_ALUCtrlD = reset ? 24'h1 : get_alu_op; // @[cu.scala 338:24]
  assign io_ALUSrcD = get_controls[22:21]; // @[cu.scala 253:33]
  assign io_RegDstD = get_controls[24:23]; // @[cu.scala 252:33]
  assign io_ImmUnsigned = get_controls[20]; // @[cu.scala 254:35]
  assign io_LinkD = 6'h0 == OpD ? 6'h9 == FunctD : _io_LinkD_T_9; // @[Mux.scala 81:58]
  assign io_HiLoWriteD = get_controls[10:9]; // @[cu.scala 259:33]
  assign io_HiLoToRegD = get_controls[8:7]; // @[cu.scala 260:34]
  assign io_CP0WriteD = get_controls[6]; // @[cu.scala 261:34]
  assign io_CP0ToRegD = get_controls[5]; // @[cu.scala 262:34]
  assign io_LoadUnsignedD = get_controls[2]; // @[cu.scala 265:38]
  assign io_MemWidthD = get_controls[1:0]; // @[cu.scala 266:32]
  assign io_MemRLD = get_controls[28:27]; // @[cu.scala 249:36]
endmodule
module dmem(
  input         io_data_ok,
  input  [31:0] io_rdata,
  input  [31:0] io_Physisc_Address,
  input  [1:0]  io_WIDTH,
  input         io_SIGN,
  output [31:0] io_RD,
  output        io_data_pending
);
  wire [1:0] ra = io_Physisc_Address[1:0]; // @[dmem.scala 39:32]
  wire [2:0] _io_RD_T_1 = {ra,io_SIGN}; // @[Cat.scala 31:58]
  wire [5:0] io_RD_lo_lo = {io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7]}; // @[Cat.scala 31:58]
  wire [11:0] io_RD_lo = {io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_RD_lo_lo}; // @[Cat.scala 31:58]
  wire [31:0] _io_RD_T_29 = {io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_RD_lo_lo,
    io_RD_lo,io_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_32 = {1'h0,io_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [5:0] io_RD_lo_lo_1 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15]}; // @[Cat.scala 31:58]
  wire [11:0] io_RD_lo_1 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_RD_lo_lo_1}
    ; // @[Cat.scala 31:58]
  wire [31:0] _io_RD_T_60 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_RD_lo_lo_1
    ,io_RD_lo_1,io_rdata[15:8]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_63 = {1'h0,io_rdata[15:8]}; // @[Cat.scala 31:58]
  wire [5:0] io_RD_lo_lo_2 = {io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23]}; // @[Cat.scala 31:58]
  wire [11:0] io_RD_lo_2 = {io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_RD_lo_lo_2}
    ; // @[Cat.scala 31:58]
  wire [31:0] _io_RD_T_91 = {io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_RD_lo_lo_2
    ,io_RD_lo_2,io_rdata[23:16]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_94 = {1'h0,io_rdata[23:16]}; // @[Cat.scala 31:58]
  wire [5:0] io_RD_lo_lo_3 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31]}; // @[Cat.scala 31:58]
  wire [11:0] io_RD_lo_3 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_RD_lo_lo_3}
    ; // @[Cat.scala 31:58]
  wire [31:0] _io_RD_T_122 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],
    io_RD_lo_lo_3,io_RD_lo_3,io_rdata[31:24]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_125 = {1'h0,io_rdata[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _io_RD_T_127 = 3'h0 == _io_RD_T_1 ? {{23'd0}, _io_RD_T_32} : _io_RD_T_29; // @[Mux.scala 81:58]
  wire [31:0] _io_RD_T_129 = 3'h3 == _io_RD_T_1 ? _io_RD_T_60 : _io_RD_T_127; // @[Mux.scala 81:58]
  wire [31:0] _io_RD_T_131 = 3'h2 == _io_RD_T_1 ? {{23'd0}, _io_RD_T_63} : _io_RD_T_129; // @[Mux.scala 81:58]
  wire [31:0] _io_RD_T_133 = 3'h5 == _io_RD_T_1 ? _io_RD_T_91 : _io_RD_T_131; // @[Mux.scala 81:58]
  wire [31:0] _io_RD_T_135 = 3'h4 == _io_RD_T_1 ? {{23'd0}, _io_RD_T_94} : _io_RD_T_133; // @[Mux.scala 81:58]
  wire [31:0] _io_RD_T_137 = 3'h7 == _io_RD_T_1 ? _io_RD_T_122 : _io_RD_T_135; // @[Mux.scala 81:58]
  wire [31:0] _io_RD_T_139 = 3'h6 == _io_RD_T_1 ? {{23'd0}, _io_RD_T_125} : _io_RD_T_137; // @[Mux.scala 81:58]
  wire [7:0] io_RD_lo_4 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],
    io_rdata[15]}; // @[Cat.scala 31:58]
  wire [31:0] _io_RD_T_160 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15]
    ,io_rdata[15],io_RD_lo_4,io_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [16:0] _io_RD_T_163 = {1'h0,io_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [7:0] io_RD_lo_5 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],
    io_rdata[31]}; // @[Cat.scala 31:58]
  wire [31:0] _io_RD_T_183 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31]
    ,io_rdata[31],io_RD_lo_5,io_rdata[31:16]}; // @[Cat.scala 31:58]
  wire [16:0] _io_RD_T_186 = {1'h0,io_rdata[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _io_RD_T_188 = 3'h1 == _io_RD_T_1 ? _io_RD_T_160 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_RD_T_190 = 3'h0 == _io_RD_T_1 ? {{15'd0}, _io_RD_T_163} : _io_RD_T_188; // @[Mux.scala 81:58]
  wire [31:0] _io_RD_T_192 = 3'h5 == _io_RD_T_1 ? _io_RD_T_183 : _io_RD_T_190; // @[Mux.scala 81:58]
  wire [31:0] _io_RD_T_194 = 3'h4 == _io_RD_T_1 ? {{15'd0}, _io_RD_T_186} : _io_RD_T_192; // @[Mux.scala 81:58]
  wire [31:0] _io_RD_T_196 = 2'h0 == io_WIDTH ? _io_RD_T_139 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_RD_T_198 = 2'h1 == io_WIDTH ? _io_RD_T_194 : _io_RD_T_196; // @[Mux.scala 81:58]
  assign io_RD = 2'h2 == io_WIDTH ? io_rdata : _io_RD_T_198; // @[Mux.scala 81:58]
  assign io_data_pending = ~io_data_ok; // @[dmem.scala 36:24]
endmodule
module dmemreq(
  input         io_en,
  input         io_MemWriteE,
  input         io_MemToRegE,
  input  [1:0]  io_MemWidthE,
  input  [31:0] io_VAddrE,
  input  [31:0] io_WriteDataE,
  input  [1:0]  io_memrl,
  output        io_req,
  output        io_wr,
  output [1:0]  io_size,
  output [31:0] io_addr,
  output [31:0] io_wdata,
  output [3:0]  io_wstrb
);
  wire [1:0] ra = io_VAddrE[1:0]; // @[dmemreq.scala 82:23]
  wire [1:0] _io_addr_T_3 = io_memrl != 2'h0 ? 2'h0 : ra; // @[dmemreq.scala 95:43]
  wire [3:0] _io_wstrb_T_1 = 2'h0 == ra ? 4'h1 : 4'hf; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_3 = 2'h1 == ra ? 4'h3 : _io_wstrb_T_1; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_5 = 2'h2 == ra ? 4'h7 : _io_wstrb_T_3; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_7 = 2'h1 == ra ? 4'he : 4'hf; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_9 = 2'h2 == ra ? 4'hc : _io_wstrb_T_7; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_11 = 2'h3 == ra ? 4'h8 : _io_wstrb_T_9; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_12 = {io_MemWidthE,ra}; // @[Cat.scala 31:58]
  wire [3:0] _io_wstrb_T_14 = io_MemWidthE == 2'h2 ? 4'hf : 4'h0; // @[dmemreq.scala 71:54]
  wire [3:0] _io_wstrb_T_16 = 4'h0 == _io_wstrb_T_12 ? 4'h1 : _io_wstrb_T_14; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_18 = 4'h1 == _io_wstrb_T_12 ? 4'h2 : _io_wstrb_T_16; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_20 = 4'h2 == _io_wstrb_T_12 ? 4'h4 : _io_wstrb_T_18; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_22 = 4'h3 == _io_wstrb_T_12 ? 4'h8 : _io_wstrb_T_20; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_24 = 4'h4 == _io_wstrb_T_12 ? 4'h3 : _io_wstrb_T_22; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_26 = 4'h6 == _io_wstrb_T_12 ? 4'hc : _io_wstrb_T_24; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_28 = 2'h2 == io_memrl ? _io_wstrb_T_5 : 4'h0; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_30 = 2'h1 == io_memrl ? _io_wstrb_T_11 : _io_wstrb_T_28; // @[Mux.scala 81:58]
  wire [31:0] _io_wdata_T_1 = {24'h0,io_WriteDataE[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _io_wdata_T_3 = {16'h0,io_WriteDataE[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _io_wdata_T_5 = {8'h0,io_WriteDataE[31:8]}; // @[Cat.scala 31:58]
  wire [31:0] _io_wdata_T_7 = 2'h0 == ra ? _io_wdata_T_1 : io_WriteDataE; // @[Mux.scala 81:58]
  wire [31:0] _io_wdata_T_9 = 2'h1 == ra ? _io_wdata_T_3 : _io_wdata_T_7; // @[Mux.scala 81:58]
  wire [31:0] _io_wdata_T_11 = 2'h2 == ra ? _io_wdata_T_5 : _io_wdata_T_9; // @[Mux.scala 81:58]
  wire [31:0] _io_wdata_T_13 = {io_WriteDataE[23:0],8'h0}; // @[Cat.scala 31:58]
  wire [31:0] _io_wdata_T_15 = {io_WriteDataE[15:0],16'h0}; // @[Cat.scala 31:58]
  wire [31:0] _io_wdata_T_17 = {io_WriteDataE[7:0],24'h0}; // @[Cat.scala 31:58]
  wire [31:0] _io_wdata_T_19 = 2'h1 == ra ? _io_wdata_T_13 : io_WriteDataE; // @[Mux.scala 81:58]
  wire [31:0] _io_wdata_T_21 = 2'h2 == ra ? _io_wdata_T_15 : _io_wdata_T_19; // @[Mux.scala 81:58]
  wire [31:0] _io_wdata_T_23 = 2'h3 == ra ? _io_wdata_T_17 : _io_wdata_T_21; // @[Mux.scala 81:58]
  wire [3:0] _io_wdata_T_24 = {ra,io_MemWidthE}; // @[Cat.scala 31:58]
  wire [31:0] _io_wdata_T_26 = {24'h0,io_WriteDataE[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_wdata_T_28 = {16'h0,io_WriteDataE[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_wdata_T_30 = {16'h0,io_WriteDataE[7:0],8'h0}; // @[Cat.scala 31:58]
  wire [31:0] _io_wdata_T_32 = {8'h0,io_WriteDataE[7:0],16'h0}; // @[Cat.scala 31:58]
  wire [31:0] _io_wdata_T_38 = 4'h0 == _io_wdata_T_24 ? _io_wdata_T_26 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_wdata_T_40 = 4'h1 == _io_wdata_T_24 ? _io_wdata_T_28 : _io_wdata_T_38; // @[Mux.scala 81:58]
  wire [31:0] _io_wdata_T_42 = 4'h2 == _io_wdata_T_24 ? io_WriteDataE : _io_wdata_T_40; // @[Mux.scala 81:58]
  wire [31:0] _io_wdata_T_44 = 4'h4 == _io_wdata_T_24 ? _io_wdata_T_30 : _io_wdata_T_42; // @[Mux.scala 81:58]
  wire [31:0] _io_wdata_T_46 = 4'h8 == _io_wdata_T_24 ? _io_wdata_T_32 : _io_wdata_T_44; // @[Mux.scala 81:58]
  wire [31:0] _io_wdata_T_48 = 4'h9 == _io_wdata_T_24 ? _io_wdata_T_15 : _io_wdata_T_46; // @[Mux.scala 81:58]
  wire [31:0] _io_wdata_T_50 = 4'hc == _io_wdata_T_24 ? _io_wdata_T_17 : _io_wdata_T_48; // @[Mux.scala 81:58]
  wire [31:0] _io_wdata_T_52 = 2'h2 == io_memrl ? _io_wdata_T_11 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_wdata_T_54 = 2'h1 == io_memrl ? _io_wdata_T_23 : _io_wdata_T_52; // @[Mux.scala 81:58]
  assign io_req = io_en & (io_MemToRegE | io_MemWriteE); // @[dmemreq.scala 98:33]
  assign io_wr = io_MemWriteE; // @[dmemreq.scala 84:17]
  assign io_size = io_MemWidthE; // @[dmemreq.scala 94:17]
  assign io_addr = {io_VAddrE[31:2],_io_addr_T_3}; // @[Cat.scala 31:58]
  assign io_wdata = 2'h0 == io_memrl ? _io_wdata_T_50 : _io_wdata_T_54; // @[Mux.scala 81:58]
  assign io_wstrb = 2'h0 == io_memrl ? _io_wstrb_T_26 : _io_wstrb_T_30; // @[Mux.scala 81:58]
endmodule
module ex2mem(
  input         clock,
  input         reset,
  input         io1_RegWriteE,
  input         io1_MemToRegE,
  input         io1_LoadUnsignedE,
  input  [1:0]  io1_MemWidthE,
  input  [1:0]  io1_HiLoWriteE,
  input         io1_CP0WriteE,
  input  [4:0]  io1_WriteCP0AddrE,
  input  [2:0]  io1_WriteCP0SelE,
  input  [31:0] io1_PCE,
  input         io1_InDelaySlotE,
  input  [1:0]  io1_MemRLE,
  input  [1:0]  io1_BranchJump_JrE,
  input  [2:0]  io1_Tlb_Control,
  input         io_en,
  input         io_clr,
  input  [4:0]  io_WriteRegE,
  input  [31:0] io_PhyAddrE,
  input  [31:0] io_HiLoOutE,
  input  [31:0] io_HiInE,
  input  [31:0] io_LoInE,
  input  [31:0] io_WriteCP0HiLoDataE,
  input  [31:0] io_BadVAddrE,
  input  [31:0] io_ExceptionTypeE,
  input  [31:0] io_RtE,
  output        io_RegWriteM,
  output        io_MemToRegM,
  output [4:0]  io_WriteRegM,
  output        io_LoadUnsignedM,
  output [1:0]  io_MemWidthM,
  output [31:0] io_PhyAddrM,
  output [1:0]  io_HiLoWriteM,
  output [31:0] io_HiLoOutM,
  output [31:0] io_HiInM,
  output [31:0] io_LoInM,
  output        io_CP0WriteM,
  output [4:0]  io_WriteCP0AddrM,
  output [2:0]  io_WriteCP0SelM,
  output [31:0] io_WriteCP0HiLoDataM,
  output [31:0] io_PCM,
  output        io_InDelaySlotM,
  output [31:0] io_BadVAddrM,
  output [31:0] io_ExceptionTypeM_Out,
  output [1:0]  io_MemRLM,
  output [31:0] io_RtM,
  output [1:0]  io_BranchJump_JrM,
  output [2:0]  io_Tlb_ControlM
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  reg  RegWrite_Reg; // @[ex2mem.scala 74:38]
  reg  MemToReg_Reg; // @[ex2mem.scala 75:38]
  reg [4:0] WriteReg_Reg; // @[ex2mem.scala 79:38]
  reg  LoadUnsigned_Reg; // @[ex2mem.scala 82:42]
  reg [1:0] MemWidth_Reg; // @[ex2mem.scala 83:38]
  reg [31:0] PhyAddr_Reg; // @[ex2mem.scala 84:37]
  reg [1:0] HiLoWrite_Reg; // @[ex2mem.scala 85:39]
  reg [31:0] HiLoOut_Reg; // @[ex2mem.scala 87:37]
  reg [31:0] HiIn_Reg; // @[ex2mem.scala 88:34]
  reg [31:0] LoIn_Reg; // @[ex2mem.scala 89:34]
  reg  CP0Write_Reg; // @[ex2mem.scala 90:38]
  reg [4:0] WriteCP0Addr_Reg; // @[ex2mem.scala 92:42]
  reg [2:0] WriteCP0Sel_Reg; // @[ex2mem.scala 93:41]
  reg [31:0] WriteCP0HiLoData_Reg; // @[ex2mem.scala 94:46]
  reg [31:0] PC_Reg; // @[ex2mem.scala 96:32]
  reg  InDelaySlot_Reg; // @[ex2mem.scala 97:41]
  reg [31:0] BadVAddr_Reg; // @[ex2mem.scala 98:38]
  reg [31:0] ExceptionType_Reg; // @[ex2mem.scala 99:41]
  reg [1:0] MemRLM_Reg; // @[ex2mem.scala 100:40]
  reg [31:0] RtM_Reg; // @[ex2mem.scala 101:32]
  reg [1:0] BranchJump_JrM_Reg; // @[ex2mem.scala 102:43]
  reg [2:0] Tlb_Control_Reg; // @[ex2mem.scala 103:43]
  assign io_RegWriteM = RegWrite_Reg; // @[ex2mem.scala 138:30]
  assign io_MemToRegM = MemToReg_Reg; // @[ex2mem.scala 139:30]
  assign io_WriteRegM = WriteReg_Reg; // @[ex2mem.scala 143:30]
  assign io_LoadUnsignedM = LoadUnsigned_Reg; // @[ex2mem.scala 146:30]
  assign io_MemWidthM = MemWidth_Reg; // @[ex2mem.scala 147:30]
  assign io_PhyAddrM = PhyAddr_Reg; // @[ex2mem.scala 148:30]
  assign io_HiLoWriteM = HiLoWrite_Reg; // @[ex2mem.scala 149:30]
  assign io_HiLoOutM = HiLoOut_Reg; // @[ex2mem.scala 151:30]
  assign io_HiInM = HiIn_Reg; // @[ex2mem.scala 152:30]
  assign io_LoInM = LoIn_Reg; // @[ex2mem.scala 153:30]
  assign io_CP0WriteM = CP0Write_Reg; // @[ex2mem.scala 154:30]
  assign io_WriteCP0AddrM = WriteCP0Addr_Reg; // @[ex2mem.scala 156:30]
  assign io_WriteCP0SelM = WriteCP0Sel_Reg; // @[ex2mem.scala 157:30]
  assign io_WriteCP0HiLoDataM = WriteCP0HiLoData_Reg; // @[ex2mem.scala 158:30]
  assign io_PCM = PC_Reg; // @[ex2mem.scala 160:30]
  assign io_InDelaySlotM = InDelaySlot_Reg; // @[ex2mem.scala 161:30]
  assign io_BadVAddrM = BadVAddr_Reg; // @[ex2mem.scala 162:30]
  assign io_ExceptionTypeM_Out = ExceptionType_Reg; // @[ex2mem.scala 163:30]
  assign io_MemRLM = MemRLM_Reg; // @[ex2mem.scala 164:30]
  assign io_RtM = RtM_Reg; // @[ex2mem.scala 165:30]
  assign io_BranchJump_JrM = BranchJump_JrM_Reg; // @[ex2mem.scala 166:30]
  assign io_Tlb_ControlM = Tlb_Control_Reg; // @[ex2mem.scala 167:30]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 105:38]
      RegWrite_Reg <= 1'h0;
    end else if (io_clr) begin // @[ex2mem.scala 105:61]
      RegWrite_Reg <= 1'h0;
    end else if (io_en) begin
      RegWrite_Reg <= io1_RegWriteE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 130:38]
      MemToReg_Reg <= 1'h0;
    end else if (io_clr) begin // @[ex2mem.scala 130:61]
      MemToReg_Reg <= 1'h0;
    end else if (io_en) begin
      MemToReg_Reg <= io1_MemToRegE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 109:38]
      WriteReg_Reg <= 5'h0;
    end else if (io_clr) begin // @[ex2mem.scala 109:61]
      WriteReg_Reg <= 5'h0;
    end else if (io_en) begin
      WriteReg_Reg <= io_WriteRegE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 112:38]
      LoadUnsigned_Reg <= 1'h0;
    end else if (io_clr) begin // @[ex2mem.scala 112:61]
      LoadUnsigned_Reg <= 1'h0;
    end else if (io_en) begin
      LoadUnsigned_Reg <= io1_LoadUnsignedE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 113:38]
      MemWidth_Reg <= 2'h0;
    end else if (io_clr) begin // @[ex2mem.scala 113:61]
      MemWidth_Reg <= 2'h0;
    end else if (io_en) begin
      MemWidth_Reg <= io1_MemWidthE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 114:38]
      PhyAddr_Reg <= 32'h0;
    end else if (io_clr) begin // @[ex2mem.scala 114:61]
      PhyAddr_Reg <= 32'h0;
    end else if (io_en) begin
      PhyAddr_Reg <= io_PhyAddrE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 115:38]
      HiLoWrite_Reg <= 2'h0;
    end else if (io_clr) begin // @[ex2mem.scala 115:61]
      HiLoWrite_Reg <= 2'h0;
    end else if (io_en) begin
      HiLoWrite_Reg <= io1_HiLoWriteE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 117:38]
      HiLoOut_Reg <= 32'h0;
    end else if (io_clr) begin // @[ex2mem.scala 117:61]
      HiLoOut_Reg <= 32'h0;
    end else if (io_en) begin
      HiLoOut_Reg <= io_HiLoOutE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 118:38]
      HiIn_Reg <= 32'h0;
    end else if (io_clr) begin // @[ex2mem.scala 118:61]
      HiIn_Reg <= 32'h0;
    end else if (io_en) begin
      HiIn_Reg <= io_HiInE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 119:38]
      LoIn_Reg <= 32'h0;
    end else if (io_clr) begin // @[ex2mem.scala 119:61]
      LoIn_Reg <= 32'h0;
    end else if (io_en) begin
      LoIn_Reg <= io_LoInE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 120:38]
      CP0Write_Reg <= 1'h0;
    end else if (io_clr) begin // @[ex2mem.scala 120:61]
      CP0Write_Reg <= 1'h0;
    end else if (io_en) begin
      CP0Write_Reg <= io1_CP0WriteE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 122:38]
      WriteCP0Addr_Reg <= 5'h0;
    end else if (io_clr) begin // @[ex2mem.scala 122:61]
      WriteCP0Addr_Reg <= 5'h0;
    end else if (io_en) begin
      WriteCP0Addr_Reg <= io1_WriteCP0AddrE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 123:38]
      WriteCP0Sel_Reg <= 3'h0;
    end else if (io_clr) begin // @[ex2mem.scala 123:61]
      WriteCP0Sel_Reg <= 3'h0;
    end else if (io_en) begin
      WriteCP0Sel_Reg <= io1_WriteCP0SelE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 124:38]
      WriteCP0HiLoData_Reg <= 32'h0;
    end else if (io_clr) begin // @[ex2mem.scala 124:61]
      WriteCP0HiLoData_Reg <= 32'h0;
    end else if (io_en) begin
      WriteCP0HiLoData_Reg <= io_WriteCP0HiLoDataE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 126:38]
      PC_Reg <= 32'h0;
    end else if (io_clr) begin // @[ex2mem.scala 126:61]
      PC_Reg <= 32'h0;
    end else if (io_en) begin
      PC_Reg <= io1_PCE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 127:38]
      InDelaySlot_Reg <= 1'h0;
    end else if (io_clr) begin // @[ex2mem.scala 127:61]
      InDelaySlot_Reg <= 1'h0;
    end else if (io_en) begin
      InDelaySlot_Reg <= io1_InDelaySlotE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 128:38]
      BadVAddr_Reg <= 32'h0;
    end else if (io_clr) begin // @[ex2mem.scala 128:61]
      BadVAddr_Reg <= 32'h0;
    end else if (io_en) begin
      BadVAddr_Reg <= io_BadVAddrE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 129:38]
      ExceptionType_Reg <= 32'h0;
    end else if (io_clr) begin // @[ex2mem.scala 129:61]
      ExceptionType_Reg <= 32'h0;
    end else if (io_en) begin
      ExceptionType_Reg <= io_ExceptionTypeE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 131:38]
      MemRLM_Reg <= 2'h0;
    end else if (io_clr) begin // @[ex2mem.scala 131:61]
      MemRLM_Reg <= 2'h0;
    end else if (io_en) begin
      MemRLM_Reg <= io1_MemRLE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 132:38]
      RtM_Reg <= 32'h0;
    end else if (io_clr) begin // @[ex2mem.scala 132:60]
      RtM_Reg <= 32'h0;
    end else if (io_en) begin
      RtM_Reg <= io_RtE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 133:38]
      BranchJump_JrM_Reg <= 2'h0;
    end else if (io_clr) begin // @[ex2mem.scala 133:60]
      BranchJump_JrM_Reg <= 2'h0;
    end else if (io_en) begin
      BranchJump_JrM_Reg <= io1_BranchJump_JrE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 134:38]
      Tlb_Control_Reg <= 3'h0;
    end else if (io_clr) begin // @[ex2mem.scala 134:61]
      Tlb_Control_Reg <= 3'h0;
    end else if (io_en) begin
      Tlb_Control_Reg <= io1_Tlb_Control;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  RegWrite_Reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  MemToReg_Reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  WriteReg_Reg = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  LoadUnsigned_Reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  MemWidth_Reg = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  PhyAddr_Reg = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  HiLoWrite_Reg = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  HiLoOut_Reg = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  HiIn_Reg = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  LoIn_Reg = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  CP0Write_Reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  WriteCP0Addr_Reg = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  WriteCP0Sel_Reg = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  WriteCP0HiLoData_Reg = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  PC_Reg = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  InDelaySlot_Reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  BadVAddr_Reg = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  ExceptionType_Reg = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  MemRLM_Reg = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  RtM_Reg = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  BranchJump_JrM_Reg = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  Tlb_Control_Reg = _RAND_21[2:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    RegWrite_Reg = 1'h0;
  end
  if (reset) begin
    MemToReg_Reg = 1'h0;
  end
  if (reset) begin
    WriteReg_Reg = 5'h0;
  end
  if (reset) begin
    LoadUnsigned_Reg = 1'h0;
  end
  if (reset) begin
    MemWidth_Reg = 2'h0;
  end
  if (reset) begin
    PhyAddr_Reg = 32'h0;
  end
  if (reset) begin
    HiLoWrite_Reg = 2'h0;
  end
  if (reset) begin
    HiLoOut_Reg = 32'h0;
  end
  if (reset) begin
    HiIn_Reg = 32'h0;
  end
  if (reset) begin
    LoIn_Reg = 32'h0;
  end
  if (reset) begin
    CP0Write_Reg = 1'h0;
  end
  if (reset) begin
    WriteCP0Addr_Reg = 5'h0;
  end
  if (reset) begin
    WriteCP0Sel_Reg = 3'h0;
  end
  if (reset) begin
    WriteCP0HiLoData_Reg = 32'h0;
  end
  if (reset) begin
    PC_Reg = 32'h0;
  end
  if (reset) begin
    InDelaySlot_Reg = 1'h0;
  end
  if (reset) begin
    BadVAddr_Reg = 32'h0;
  end
  if (reset) begin
    ExceptionType_Reg = 32'h0;
  end
  if (reset) begin
    MemRLM_Reg = 2'h0;
  end
  if (reset) begin
    RtM_Reg = 32'h0;
  end
  if (reset) begin
    BranchJump_JrM_Reg = 2'h0;
  end
  if (reset) begin
    Tlb_Control_Reg = 3'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module hilo(
  input         clock,
  input         reset,
  input  [1:0]  io_we,
  input  [31:0] io_hi_i,
  input  [31:0] io_lo_i,
  output [31:0] io_hi_o,
  output [31:0] io_lo_o
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] hi_o_Reg; // @[hilo.scala 20:30]
  reg [31:0] lo_o_Reg; // @[hilo.scala 21:30]
  assign io_hi_o = hi_o_Reg; // @[hilo.scala 22:17]
  assign io_lo_o = lo_o_Reg; // @[hilo.scala 23:17]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hilo.scala 26:20]
      hi_o_Reg <= 32'h0;
    end else if (io_we[1]) begin
      hi_o_Reg <= io_hi_i;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hilo.scala 25:20]
      lo_o_Reg <= 32'h0;
    end else if (io_we[0]) begin
      lo_o_Reg <= io_lo_i;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hi_o_Reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  lo_o_Reg = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    hi_o_Reg = 32'h0;
  end
  if (reset) begin
    lo_o_Reg = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module id2ex(
  input         clock,
  input         reset,
  input         io1_RegWriteD,
  input         io1_MemToRegD,
  input         io1_MemWriteD,
  input  [23:0] io1_ALUCtrlD,
  input  [1:0]  io1_ALUSrcD,
  input  [1:0]  io1_RegDstD,
  input         io1_LinkD,
  input  [1:0]  io1_HiLoWriteD,
  input  [1:0]  io1_HiLoToRegD,
  input         io1_CP0WriteD,
  input         io1_CP0ToRegD,
  input         io1_LoadUnsignedD,
  input  [1:0]  io1_MemWidthD,
  input  [1:0]  io1_MemRLD,
  output        io2_RegWriteE,
  output        io2_MemToRegE,
  output        io2_MemWriteE,
  output [23:0] io2_ALUCtrlE,
  output [1:0]  io2_ALUSrcE,
  output [1:0]  io2_RegDstE,
  output        io2_LinkE,
  output [31:0] io2_PCPlus8E,
  output        io2_LoadUnsignedE,
  output [1:0]  io2_MemWidthE,
  output [1:0]  io2_HiLoWriteE,
  output [1:0]  io2_HiLoToRegE,
  output        io2_CP0WriteE,
  output [4:0]  io2_WriteCP0AddrE,
  output [2:0]  io2_WriteCP0SelE,
  output [4:0]  io2_ReadCP0AddrE,
  output [2:0]  io2_ReadCP0SelE,
  output [31:0] io2_PCE,
  output        io2_InDelaySlotE,
  output [1:0]  io2_MemRLE,
  output [1:0]  io2_BranchJump_JrE,
  output [2:0]  io2_Tlb_Control,
  input         io_en,
  input         io_clr,
  output        io_CP0ToRegE_Out,
  input  [31:0] io_RD1D,
  input  [31:0] io_RD2D,
  input  [4:0]  io_RsD,
  input  [4:0]  io_RtD,
  input  [4:0]  io_RdD,
  input  [31:0] io_ImmD,
  input  [31:0] io_PCPlus8D,
  input  [4:0]  io_WriteCP0AddrD,
  input  [2:0]  io_WriteCP0SelD,
  input  [4:0]  io_ReadCP0AddrD,
  input  [2:0]  io_ReadCP0SelD,
  input  [31:0] io_PCD,
  input         io_InDelaySlotD,
  input  [31:0] io_ExceptionTypeD,
  input  [1:0]  io_BranchJump_JrD,
  input  [31:0] io_BadVaddrD,
  input  [2:0]  io_Tlb_Control,
  output [31:0] io_RD1E,
  output [31:0] io_RD2E,
  output [4:0]  io_RsE,
  output [4:0]  io_RtE,
  output [4:0]  io_RdE,
  output [31:0] io_ImmE,
  output [31:0] io_BadVaddrE,
  output [31:0] io_ExceptionTypeE_Out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg  RegWriteE_Reg; // @[id2ex.scala 118:35]
  reg  MemToRegE_Reg; // @[id2ex.scala 119:35]
  reg  MemWriteE_Reg; // @[id2ex.scala 120:35]
  reg [23:0] ALUCtrlE_Reg; // @[id2ex.scala 121:34]
  reg [1:0] ALUSrcE_Reg; // @[id2ex.scala 122:33]
  reg [1:0] RegDstE_Reg; // @[id2ex.scala 123:33]
  reg [31:0] RD1E_Reg; // @[id2ex.scala 124:30]
  reg [31:0] RD2E_Reg; // @[id2ex.scala 125:30]
  reg [4:0] RsE_Reg; // @[id2ex.scala 126:29]
  reg [4:0] RtE_Reg; // @[id2ex.scala 127:29]
  reg [4:0] RdE_Reg; // @[id2ex.scala 128:29]
  reg [31:0] ImmE_Reg; // @[id2ex.scala 129:30]
  reg  LinkE_Reg; // @[id2ex.scala 130:31]
  reg [31:0] PCPlus8E_Reg; // @[id2ex.scala 131:34]
  reg  LoadUnsignedE_Reg; // @[id2ex.scala 132:39]
  reg [1:0] MemWidthE_Reg; // @[id2ex.scala 133:35]
  reg [1:0] HiLoWriteE_Reg; // @[id2ex.scala 134:36]
  reg [1:0] HiLoToRegE_Reg; // @[id2ex.scala 135:36]
  reg  CP0WriteE_Reg; // @[id2ex.scala 136:35]
  reg  CP0ToRegE_Reg; // @[id2ex.scala 137:35]
  reg [4:0] WriteCP0AddrE_Reg; // @[id2ex.scala 138:39]
  reg [2:0] WriteCP0SelE_Reg; // @[id2ex.scala 139:38]
  reg [4:0] ReadCP0AddrE_Reg; // @[id2ex.scala 140:38]
  reg [2:0] ReadCP0SelE_Reg; // @[id2ex.scala 141:37]
  reg [31:0] PCE_Reg; // @[id2ex.scala 142:29]
  reg  InDelaySlotE_Reg; // @[id2ex.scala 143:38]
  reg [31:0] ExceptionTypeE_Reg; // @[id2ex.scala 144:40]
  reg [1:0] MemRLE_Reg; // @[id2ex.scala 145:38]
  reg [1:0] BranchJump_JrE_Reg; // @[id2ex.scala 146:40]
  reg [31:0] BadVaddrE_Reg; // @[id2ex.scala 147:35]
  reg [2:0] Tlb_Control_Reg; // @[id2ex.scala 148:39]
  assign io2_RegWriteE = RegWriteE_Reg; // @[id2ex.scala 183:33]
  assign io2_MemToRegE = MemToRegE_Reg; // @[id2ex.scala 184:33]
  assign io2_MemWriteE = MemWriteE_Reg; // @[id2ex.scala 185:23]
  assign io2_ALUCtrlE = ALUCtrlE_Reg; // @[id2ex.scala 186:23]
  assign io2_ALUSrcE = ALUSrcE_Reg; // @[id2ex.scala 187:23]
  assign io2_RegDstE = RegDstE_Reg; // @[id2ex.scala 188:23]
  assign io2_LinkE = LinkE_Reg; // @[id2ex.scala 195:23]
  assign io2_PCPlus8E = PCPlus8E_Reg; // @[id2ex.scala 196:23]
  assign io2_LoadUnsignedE = LoadUnsignedE_Reg; // @[id2ex.scala 197:23]
  assign io2_MemWidthE = MemWidthE_Reg; // @[id2ex.scala 198:23]
  assign io2_HiLoWriteE = HiLoWriteE_Reg; // @[id2ex.scala 199:23]
  assign io2_HiLoToRegE = HiLoToRegE_Reg; // @[id2ex.scala 200:23]
  assign io2_CP0WriteE = CP0WriteE_Reg; // @[id2ex.scala 201:23]
  assign io2_WriteCP0AddrE = WriteCP0AddrE_Reg; // @[id2ex.scala 203:23]
  assign io2_WriteCP0SelE = WriteCP0SelE_Reg; // @[id2ex.scala 204:23]
  assign io2_ReadCP0AddrE = ReadCP0AddrE_Reg; // @[id2ex.scala 205:23]
  assign io2_ReadCP0SelE = ReadCP0SelE_Reg; // @[id2ex.scala 206:23]
  assign io2_PCE = PCE_Reg; // @[id2ex.scala 207:23]
  assign io2_InDelaySlotE = InDelaySlotE_Reg; // @[id2ex.scala 208:23]
  assign io2_MemRLE = MemRLE_Reg; // @[id2ex.scala 209:23]
  assign io2_BranchJump_JrE = BranchJump_JrE_Reg; // @[id2ex.scala 211:24]
  assign io2_Tlb_Control = Tlb_Control_Reg; // @[id2ex.scala 213:23]
  assign io_CP0ToRegE_Out = CP0ToRegE_Reg; // @[id2ex.scala 202:26]
  assign io_RD1E = RD1E_Reg; // @[id2ex.scala 189:22]
  assign io_RD2E = RD2E_Reg; // @[id2ex.scala 190:22]
  assign io_RsE = RsE_Reg; // @[id2ex.scala 191:22]
  assign io_RtE = RtE_Reg; // @[id2ex.scala 192:22]
  assign io_RdE = RdE_Reg; // @[id2ex.scala 193:22]
  assign io_ImmE = ImmE_Reg; // @[id2ex.scala 194:22]
  assign io_BadVaddrE = BadVaddrE_Reg; // @[id2ex.scala 212:23]
  assign io_ExceptionTypeE_Out = ExceptionTypeE_Reg; // @[id2ex.scala 210:26]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 151:42]
      RegWriteE_Reg <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 151:64]
      RegWriteE_Reg <= 1'h0;
    end else if (io_en) begin
      RegWriteE_Reg <= io1_RegWriteD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 152:42]
      MemToRegE_Reg <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 152:64]
      MemToRegE_Reg <= 1'h0;
    end else if (io_en) begin
      MemToRegE_Reg <= io1_MemToRegD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 153:42]
      MemWriteE_Reg <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 153:64]
      MemWriteE_Reg <= 1'h0;
    end else if (io_en) begin
      MemWriteE_Reg <= io1_MemWriteD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 154:42]
      ALUCtrlE_Reg <= 24'h0;
    end else if (io_clr) begin // @[id2ex.scala 154:64]
      ALUCtrlE_Reg <= 24'h0;
    end else if (io_en) begin
      ALUCtrlE_Reg <= io1_ALUCtrlD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 155:42]
      ALUSrcE_Reg <= 2'h0;
    end else if (io_clr) begin // @[id2ex.scala 155:64]
      ALUSrcE_Reg <= 2'h0;
    end else if (io_en) begin
      ALUSrcE_Reg <= io1_ALUSrcD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 156:42]
      RegDstE_Reg <= 2'h0;
    end else if (io_clr) begin // @[id2ex.scala 156:64]
      RegDstE_Reg <= 2'h0;
    end else if (io_en) begin
      RegDstE_Reg <= io1_RegDstD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 157:42]
      RD1E_Reg <= 32'h0;
    end else if (io_clr) begin // @[id2ex.scala 157:64]
      RD1E_Reg <= 32'h0;
    end else if (io_en) begin
      RD1E_Reg <= io_RD1D;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 158:42]
      RD2E_Reg <= 32'h0;
    end else if (io_clr) begin // @[id2ex.scala 158:64]
      RD2E_Reg <= 32'h0;
    end else if (io_en) begin
      RD2E_Reg <= io_RD2D;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 159:42]
      RsE_Reg <= 5'h0;
    end else if (io_clr) begin // @[id2ex.scala 159:64]
      RsE_Reg <= 5'h0;
    end else if (io_en) begin
      RsE_Reg <= io_RsD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 160:42]
      RtE_Reg <= 5'h0;
    end else if (io_clr) begin // @[id2ex.scala 160:64]
      RtE_Reg <= 5'h0;
    end else if (io_en) begin
      RtE_Reg <= io_RtD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 161:42]
      RdE_Reg <= 5'h0;
    end else if (io_clr) begin // @[id2ex.scala 161:64]
      RdE_Reg <= 5'h0;
    end else if (io_en) begin
      RdE_Reg <= io_RdD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 162:42]
      ImmE_Reg <= 32'h0;
    end else if (io_clr) begin // @[id2ex.scala 162:64]
      ImmE_Reg <= 32'h0;
    end else if (io_en) begin
      ImmE_Reg <= io_ImmD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 163:42]
      LinkE_Reg <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 163:64]
      LinkE_Reg <= 1'h0;
    end else if (io_en) begin
      LinkE_Reg <= io1_LinkD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 164:42]
      PCPlus8E_Reg <= 32'h0;
    end else if (io_clr) begin // @[id2ex.scala 164:64]
      PCPlus8E_Reg <= 32'h0;
    end else if (io_en) begin
      PCPlus8E_Reg <= io_PCPlus8D;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 165:42]
      LoadUnsignedE_Reg <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 165:64]
      LoadUnsignedE_Reg <= 1'h0;
    end else if (io_en) begin
      LoadUnsignedE_Reg <= io1_LoadUnsignedD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 166:42]
      MemWidthE_Reg <= 2'h0;
    end else if (io_clr) begin // @[id2ex.scala 166:64]
      MemWidthE_Reg <= 2'h0;
    end else if (io_en) begin
      MemWidthE_Reg <= io1_MemWidthD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 167:42]
      HiLoWriteE_Reg <= 2'h0;
    end else if (io_clr) begin // @[id2ex.scala 167:64]
      HiLoWriteE_Reg <= 2'h0;
    end else if (io_en) begin
      HiLoWriteE_Reg <= io1_HiLoWriteD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 168:42]
      HiLoToRegE_Reg <= 2'h0;
    end else if (io_clr) begin // @[id2ex.scala 168:64]
      HiLoToRegE_Reg <= 2'h0;
    end else if (io_en) begin
      HiLoToRegE_Reg <= io1_HiLoToRegD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 169:42]
      CP0WriteE_Reg <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 169:64]
      CP0WriteE_Reg <= 1'h0;
    end else if (io_en) begin
      CP0WriteE_Reg <= io1_CP0WriteD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 170:42]
      CP0ToRegE_Reg <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 170:64]
      CP0ToRegE_Reg <= 1'h0;
    end else if (io_en) begin
      CP0ToRegE_Reg <= io1_CP0ToRegD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 171:42]
      WriteCP0AddrE_Reg <= 5'h0;
    end else if (io_clr) begin // @[id2ex.scala 171:64]
      WriteCP0AddrE_Reg <= 5'h0;
    end else if (io_en) begin
      WriteCP0AddrE_Reg <= io_WriteCP0AddrD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 172:42]
      WriteCP0SelE_Reg <= 3'h0;
    end else if (io_clr) begin // @[id2ex.scala 172:64]
      WriteCP0SelE_Reg <= 3'h0;
    end else if (io_en) begin
      WriteCP0SelE_Reg <= io_WriteCP0SelD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 173:42]
      ReadCP0AddrE_Reg <= 5'h0;
    end else if (io_clr) begin // @[id2ex.scala 173:64]
      ReadCP0AddrE_Reg <= 5'h0;
    end else if (io_en) begin
      ReadCP0AddrE_Reg <= io_ReadCP0AddrD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 174:42]
      ReadCP0SelE_Reg <= 3'h0;
    end else if (io_clr) begin // @[id2ex.scala 174:64]
      ReadCP0SelE_Reg <= 3'h0;
    end else if (io_en) begin
      ReadCP0SelE_Reg <= io_ReadCP0SelD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 175:42]
      PCE_Reg <= 32'h0;
    end else if (io_clr) begin // @[id2ex.scala 175:64]
      PCE_Reg <= 32'h0;
    end else if (io_en) begin
      PCE_Reg <= io_PCD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 176:42]
      InDelaySlotE_Reg <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 176:64]
      InDelaySlotE_Reg <= 1'h0;
    end else if (io_en) begin
      InDelaySlotE_Reg <= io_InDelaySlotD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 177:42]
      ExceptionTypeE_Reg <= 32'h0;
    end else if (io_clr) begin // @[id2ex.scala 177:64]
      ExceptionTypeE_Reg <= 32'h0;
    end else if (io_en) begin
      ExceptionTypeE_Reg <= io_ExceptionTypeD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 178:42]
      MemRLE_Reg <= 2'h0;
    end else if (io_clr) begin // @[id2ex.scala 178:64]
      MemRLE_Reg <= 2'h0;
    end else if (io_en) begin
      MemRLE_Reg <= io1_MemRLD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 179:42]
      BranchJump_JrE_Reg <= 2'h0;
    end else if (io_clr) begin // @[id2ex.scala 179:64]
      BranchJump_JrE_Reg <= 2'h0;
    end else if (io_en) begin
      BranchJump_JrE_Reg <= io_BranchJump_JrD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 180:42]
      BadVaddrE_Reg <= 32'h0;
    end else if (io_clr) begin // @[id2ex.scala 180:64]
      BadVaddrE_Reg <= 32'h0;
    end else if (io_en) begin
      BadVaddrE_Reg <= io_BadVaddrD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 181:42]
      Tlb_Control_Reg <= 3'h0;
    end else if (io_clr) begin // @[id2ex.scala 181:64]
      Tlb_Control_Reg <= 3'h0;
    end else if (io_en) begin
      Tlb_Control_Reg <= io_Tlb_Control;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  RegWriteE_Reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  MemToRegE_Reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  MemWriteE_Reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ALUCtrlE_Reg = _RAND_3[23:0];
  _RAND_4 = {1{`RANDOM}};
  ALUSrcE_Reg = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  RegDstE_Reg = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  RD1E_Reg = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  RD2E_Reg = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  RsE_Reg = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  RtE_Reg = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  RdE_Reg = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  ImmE_Reg = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  LinkE_Reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  PCPlus8E_Reg = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  LoadUnsignedE_Reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  MemWidthE_Reg = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  HiLoWriteE_Reg = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  HiLoToRegE_Reg = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  CP0WriteE_Reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  CP0ToRegE_Reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  WriteCP0AddrE_Reg = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  WriteCP0SelE_Reg = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  ReadCP0AddrE_Reg = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  ReadCP0SelE_Reg = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  PCE_Reg = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  InDelaySlotE_Reg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  ExceptionTypeE_Reg = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  MemRLE_Reg = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  BranchJump_JrE_Reg = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  BadVaddrE_Reg = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  Tlb_Control_Reg = _RAND_30[2:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    RegWriteE_Reg = 1'h0;
  end
  if (reset) begin
    MemToRegE_Reg = 1'h0;
  end
  if (reset) begin
    MemWriteE_Reg = 1'h0;
  end
  if (reset) begin
    ALUCtrlE_Reg = 24'h0;
  end
  if (reset) begin
    ALUSrcE_Reg = 2'h0;
  end
  if (reset) begin
    RegDstE_Reg = 2'h0;
  end
  if (reset) begin
    RD1E_Reg = 32'h0;
  end
  if (reset) begin
    RD2E_Reg = 32'h0;
  end
  if (reset) begin
    RsE_Reg = 5'h0;
  end
  if (reset) begin
    RtE_Reg = 5'h0;
  end
  if (reset) begin
    RdE_Reg = 5'h0;
  end
  if (reset) begin
    ImmE_Reg = 32'h0;
  end
  if (reset) begin
    LinkE_Reg = 1'h0;
  end
  if (reset) begin
    PCPlus8E_Reg = 32'h0;
  end
  if (reset) begin
    LoadUnsignedE_Reg = 1'h0;
  end
  if (reset) begin
    MemWidthE_Reg = 2'h0;
  end
  if (reset) begin
    HiLoWriteE_Reg = 2'h0;
  end
  if (reset) begin
    HiLoToRegE_Reg = 2'h0;
  end
  if (reset) begin
    CP0WriteE_Reg = 1'h0;
  end
  if (reset) begin
    CP0ToRegE_Reg = 1'h0;
  end
  if (reset) begin
    WriteCP0AddrE_Reg = 5'h0;
  end
  if (reset) begin
    WriteCP0SelE_Reg = 3'h0;
  end
  if (reset) begin
    ReadCP0AddrE_Reg = 5'h0;
  end
  if (reset) begin
    ReadCP0SelE_Reg = 3'h0;
  end
  if (reset) begin
    PCE_Reg = 32'h0;
  end
  if (reset) begin
    InDelaySlotE_Reg = 1'h0;
  end
  if (reset) begin
    ExceptionTypeE_Reg = 32'h0;
  end
  if (reset) begin
    MemRLE_Reg = 2'h0;
  end
  if (reset) begin
    BranchJump_JrE_Reg = 2'h0;
  end
  if (reset) begin
    BadVaddrE_Reg = 32'h0;
  end
  if (reset) begin
    Tlb_Control_Reg = 3'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module if2id(
  input         clock,
  input         reset,
  input         io_en,
  input         io_clr,
  input  [31:0] io_InstrF,
  input  [31:0] io_PCPlus4F,
  input  [31:0] io_PCPlus8F,
  input  [31:0] io_PCF,
  input  [1:0]  io_ExceptionTypeF,
  input         io_NextDelaySlotD,
  output [31:0] io_InstrD,
  output [31:0] io_PCPlus4D,
  output [31:0] io_PCPlus8D,
  output        io_InDelaySlotD,
  output [31:0] io_PCD,
  output [1:0]  io_ExceptionTypeD_Out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] InstrD_Reg; // @[if2id.scala 36:29]
  reg [31:0] PCPlus4D_Reg; // @[if2id.scala 37:31]
  reg [31:0] PCPlus8D_Reg; // @[if2id.scala 38:31]
  reg [31:0] PCD_Reg; // @[if2id.scala 39:26]
  reg [1:0] ExceptionTypeD_Reg; // @[if2id.scala 40:37]
  reg  InDelaySlotD_Reg; // @[if2id.scala 41:35]
  assign io_InstrD = InstrD_Reg; // @[if2id.scala 46:15]
  assign io_PCPlus4D = PCPlus4D_Reg; // @[if2id.scala 47:17]
  assign io_PCPlus8D = PCPlus8D_Reg; // @[if2id.scala 48:17]
  assign io_InDelaySlotD = InDelaySlotD_Reg; // @[if2id.scala 49:21]
  assign io_PCD = PCD_Reg; // @[if2id.scala 51:13]
  assign io_ExceptionTypeD_Out = ExceptionTypeD_Reg; // @[if2id.scala 50:27]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[if2id.scala 55:35]
      InstrD_Reg <= 32'h0;
    end else if (io_clr) begin // @[if2id.scala 55:57]
      InstrD_Reg <= 32'h0;
    end else if (io_en) begin
      InstrD_Reg <= io_InstrF;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[if2id.scala 56:35]
      PCPlus4D_Reg <= 32'h0;
    end else if (io_clr) begin // @[if2id.scala 56:57]
      PCPlus4D_Reg <= 32'h0;
    end else if (io_en) begin
      PCPlus4D_Reg <= io_PCPlus4F;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[if2id.scala 57:35]
      PCPlus8D_Reg <= 32'h0;
    end else if (io_clr) begin // @[if2id.scala 57:57]
      PCPlus8D_Reg <= 32'h0;
    end else if (io_en) begin
      PCPlus8D_Reg <= io_PCPlus8F;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[if2id.scala 58:39]
      PCD_Reg <= 32'h0;
    end else if (io_clr) begin // @[if2id.scala 58:61]
      PCD_Reg <= 32'h0;
    end else if (io_en) begin
      PCD_Reg <= io_PCF;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[if2id.scala 59:39]
      ExceptionTypeD_Reg <= 2'h0;
    end else if (io_clr) begin // @[if2id.scala 59:61]
      ExceptionTypeD_Reg <= 2'h0;
    end else if (io_en) begin
      ExceptionTypeD_Reg <= io_ExceptionTypeF;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[if2id.scala 60:39]
      InDelaySlotD_Reg <= 1'h0;
    end else if (io_clr) begin // @[if2id.scala 60:61]
      InDelaySlotD_Reg <= 1'h0;
    end else if (io_en) begin
      InDelaySlotD_Reg <= io_NextDelaySlotD;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  InstrD_Reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  PCPlus4D_Reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  PCPlus8D_Reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  PCD_Reg = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  ExceptionTypeD_Reg = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  InDelaySlotD_Reg = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    InstrD_Reg = 32'h0;
  end
  if (reset) begin
    PCPlus4D_Reg = 32'h0;
  end
  if (reset) begin
    PCPlus8D_Reg = 32'h0;
  end
  if (reset) begin
    PCD_Reg = 32'h0;
  end
  if (reset) begin
    ExceptionTypeD_Reg = 2'h0;
  end
  if (reset) begin
    InDelaySlotD_Reg = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module mem2wb(
  input         clock,
  input         reset,
  input         io_en,
  input         io_clr,
  input         io_RegWriteM,
  input  [31:0] io_ResultM,
  input  [4:0]  io_WriteRegM,
  input  [1:0]  io_HiLoWriteM,
  input  [31:0] io_HiInM,
  input  [31:0] io_LoInM,
  input         io_CP0WriteM,
  input  [4:0]  io_WriteCP0AddrM,
  input  [2:0]  io_WriteCP0SelM,
  input  [31:0] io_WriteCP0HiLoDataM,
  input  [31:0] io_PCM,
  input         io_InDelaySlotM,
  input  [31:0] io_BadVAddrM,
  input  [31:0] io_ExceptionTypeM,
  input  [1:0]  io_BranchJump_JrM,
  input  [2:0]  io_Tlb_ControlM,
  output        io_RegWriteW_Out,
  output [31:0] io_ResultW,
  output [4:0]  io_WriteRegW,
  output [1:0]  io_HiLoWriteW,
  output [31:0] io_HiInW,
  output [31:0] io_LoInW,
  output        io_CP0WriteW,
  output [4:0]  io_WriteCP0AddrW,
  output [2:0]  io_WriteCP0SelW,
  output [31:0] io_WriteCP0HiLoDataW,
  output [31:0] io_PCW,
  output        io_InDelaySlotW,
  output [31:0] io_BadVAddrW,
  output [31:0] io_ExceptionTypeW_Out,
  output [1:0]  io_BranchJump_JrW,
  output [2:0]  io_Tlb_ControlW
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg  RegWriteW; // @[mem2wb.scala 57:34]
  reg [31:0] ResultW; // @[mem2wb.scala 60:32]
  reg [4:0] WriteRegW; // @[mem2wb.scala 61:34]
  reg [1:0] HiLoWriteW; // @[mem2wb.scala 62:35]
  reg [31:0] HiInW; // @[mem2wb.scala 63:30]
  reg [31:0] LoInW; // @[mem2wb.scala 64:30]
  reg  CP0WriteW; // @[mem2wb.scala 65:34]
  reg [4:0] WriteCP0AddrW; // @[mem2wb.scala 66:38]
  reg [2:0] WriteCP0SelW; // @[mem2wb.scala 67:37]
  reg [31:0] WriteCP0HiLoDataW; // @[mem2wb.scala 68:42]
  reg [31:0] PCW; // @[mem2wb.scala 69:28]
  reg  InDelaySlotW; // @[mem2wb.scala 70:37]
  reg [31:0] BadVAddrW; // @[mem2wb.scala 71:34]
  reg [31:0] ExceptionTypeW; // @[mem2wb.scala 72:39]
  reg [1:0] BranchJump_JrW_Reg; // @[mem2wb.scala 74:43]
  reg [2:0] Tlb_Control_Reg; // @[mem2wb.scala 75:40]
  assign io_RegWriteW_Out = RegWriteW; // @[mem2wb.scala 78:36]
  assign io_ResultW = ResultW; // @[mem2wb.scala 81:32]
  assign io_WriteRegW = WriteRegW; // @[mem2wb.scala 82:32]
  assign io_HiLoWriteW = HiLoWriteW; // @[mem2wb.scala 83:32]
  assign io_HiInW = HiInW; // @[mem2wb.scala 84:32]
  assign io_LoInW = LoInW; // @[mem2wb.scala 85:32]
  assign io_CP0WriteW = CP0WriteW; // @[mem2wb.scala 86:32]
  assign io_WriteCP0AddrW = WriteCP0AddrW; // @[mem2wb.scala 87:32]
  assign io_WriteCP0SelW = WriteCP0SelW; // @[mem2wb.scala 88:32]
  assign io_WriteCP0HiLoDataW = WriteCP0HiLoDataW; // @[mem2wb.scala 89:32]
  assign io_PCW = PCW; // @[mem2wb.scala 90:32]
  assign io_InDelaySlotW = InDelaySlotW; // @[mem2wb.scala 91:32]
  assign io_BadVAddrW = BadVAddrW; // @[mem2wb.scala 92:32]
  assign io_ExceptionTypeW_Out = ExceptionTypeW; // @[mem2wb.scala 93:32]
  assign io_BranchJump_JrW = BranchJump_JrW_Reg; // @[mem2wb.scala 94:32]
  assign io_Tlb_ControlW = Tlb_Control_Reg; // @[mem2wb.scala 95:32]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 100:34]
      RegWriteW <= 1'h0;
    end else if (io_clr) begin // @[mem2wb.scala 100:56]
      RegWriteW <= 1'h0;
    end else if (io_en) begin
      RegWriteW <= io_RegWriteM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 103:34]
      ResultW <= 32'h0;
    end else if (io_clr) begin // @[mem2wb.scala 103:56]
      ResultW <= 32'h0;
    end else if (io_en) begin
      ResultW <= io_ResultM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 104:34]
      WriteRegW <= 5'h0;
    end else if (io_clr) begin // @[mem2wb.scala 104:56]
      WriteRegW <= 5'h0;
    end else if (io_en) begin
      WriteRegW <= io_WriteRegM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 105:34]
      HiLoWriteW <= 2'h0;
    end else if (io_clr) begin // @[mem2wb.scala 105:56]
      HiLoWriteW <= 2'h0;
    end else if (io_en) begin
      HiLoWriteW <= io_HiLoWriteM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 106:34]
      HiInW <= 32'h0;
    end else if (io_clr) begin // @[mem2wb.scala 106:56]
      HiInW <= 32'h0;
    end else if (io_en) begin
      HiInW <= io_HiInM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 107:34]
      LoInW <= 32'h0;
    end else if (io_clr) begin // @[mem2wb.scala 107:56]
      LoInW <= 32'h0;
    end else if (io_en) begin
      LoInW <= io_LoInM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 108:34]
      CP0WriteW <= 1'h0;
    end else if (io_clr) begin // @[mem2wb.scala 108:56]
      CP0WriteW <= 1'h0;
    end else if (io_en) begin
      CP0WriteW <= io_CP0WriteM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 109:34]
      WriteCP0AddrW <= 5'h0;
    end else if (io_clr) begin // @[mem2wb.scala 109:56]
      WriteCP0AddrW <= 5'h0;
    end else if (io_en) begin
      WriteCP0AddrW <= io_WriteCP0AddrM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 110:34]
      WriteCP0SelW <= 3'h0;
    end else if (io_clr) begin // @[mem2wb.scala 110:56]
      WriteCP0SelW <= 3'h0;
    end else if (io_en) begin
      WriteCP0SelW <= io_WriteCP0SelM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 111:34]
      WriteCP0HiLoDataW <= 32'h0;
    end else if (io_clr) begin // @[mem2wb.scala 111:56]
      WriteCP0HiLoDataW <= 32'h0;
    end else if (io_en) begin
      WriteCP0HiLoDataW <= io_WriteCP0HiLoDataM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 112:34]
      PCW <= 32'h0;
    end else if (io_clr) begin // @[mem2wb.scala 112:56]
      PCW <= 32'h0;
    end else if (io_en) begin
      PCW <= io_PCM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 113:34]
      InDelaySlotW <= 1'h0;
    end else if (io_clr) begin // @[mem2wb.scala 113:56]
      InDelaySlotW <= 1'h0;
    end else if (io_en) begin
      InDelaySlotW <= io_InDelaySlotM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 114:34]
      BadVAddrW <= 32'h0;
    end else if (io_clr) begin // @[mem2wb.scala 114:56]
      BadVAddrW <= 32'h0;
    end else if (io_en) begin
      BadVAddrW <= io_BadVAddrM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 115:34]
      ExceptionTypeW <= 32'h0;
    end else if (io_clr) begin // @[mem2wb.scala 115:56]
      ExceptionTypeW <= 32'h0;
    end else if (io_en) begin
      ExceptionTypeW <= io_ExceptionTypeM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 116:49]
      BranchJump_JrW_Reg <= 2'h0;
    end else if (io_clr) begin // @[mem2wb.scala 116:71]
      BranchJump_JrW_Reg <= 2'h0;
    end else if (io_en) begin
      BranchJump_JrW_Reg <= io_BranchJump_JrM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 117:34]
      Tlb_Control_Reg <= 3'h0;
    end else if (io_clr) begin // @[mem2wb.scala 117:56]
      Tlb_Control_Reg <= 3'h0;
    end else if (io_en) begin
      Tlb_Control_Reg <= io_Tlb_ControlM;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  RegWriteW = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ResultW = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  WriteRegW = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  HiLoWriteW = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  HiInW = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  LoInW = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  CP0WriteW = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  WriteCP0AddrW = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  WriteCP0SelW = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  WriteCP0HiLoDataW = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  PCW = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  InDelaySlotW = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  BadVAddrW = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  ExceptionTypeW = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  BranchJump_JrW_Reg = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  Tlb_Control_Reg = _RAND_15[2:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    RegWriteW = 1'h0;
  end
  if (reset) begin
    ResultW = 32'h0;
  end
  if (reset) begin
    WriteRegW = 5'h0;
  end
  if (reset) begin
    HiLoWriteW = 2'h0;
  end
  if (reset) begin
    HiInW = 32'h0;
  end
  if (reset) begin
    LoInW = 32'h0;
  end
  if (reset) begin
    CP0WriteW = 1'h0;
  end
  if (reset) begin
    WriteCP0AddrW = 5'h0;
  end
  if (reset) begin
    WriteCP0SelW = 3'h0;
  end
  if (reset) begin
    WriteCP0HiLoDataW = 32'h0;
  end
  if (reset) begin
    PCW = 32'h0;
  end
  if (reset) begin
    InDelaySlotW = 1'h0;
  end
  if (reset) begin
    BadVAddrW = 32'h0;
  end
  if (reset) begin
    ExceptionTypeW = 32'h0;
  end
  if (reset) begin
    BranchJump_JrW_Reg = 2'h0;
  end
  if (reset) begin
    Tlb_Control_Reg = 3'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module addr_cal(
  input  [31:0] io_d_vaddr,
  input  [1:0]  io_d_width,
  input  [1:0]  io_d_memrl,
  output [31:0] io_d_paddr,
  output        io_d_cached,
  output        io_d_unaligned
);
  wire [2:0] _io_d_unaligned_T_3 = {io_d_width,io_d_vaddr[0]}; // @[Cat.scala 31:58]
  wire  _io_d_unaligned_T_4 = _io_d_unaligned_T_3 == 3'h2; // @[macros.scala 417:27]
  wire [3:0] _io_d_unaligned_T_5 = {io_d_width,io_d_vaddr[1:0]}; // @[Cat.scala 31:58]
  wire  _io_d_unaligned_T_6 = _io_d_unaligned_T_5 == 4'h8; // @[macros.scala 418:24]
  wire  _io_d_unaligned_T_7 = io_d_width == 2'h0; // @[macros.scala 419:16]
  wire  _io_d_unaligned_T_8 = _io_d_unaligned_T_7 ? 1'h0 : 1'h1; // @[Mux.scala 101:16]
  wire  _io_d_unaligned_T_9 = _io_d_unaligned_T_6 ? 1'h0 : _io_d_unaligned_T_8; // @[Mux.scala 101:16]
  wire  _io_d_unaligned_T_10 = _io_d_unaligned_T_4 ? 1'h0 : _io_d_unaligned_T_9; // @[Mux.scala 101:16]
  assign io_d_paddr = io_d_vaddr; // @[addr_cal.scala 24:16]
  assign io_d_cached = io_d_vaddr[31:29] == 3'h4; // @[macros.scala 420:55]
  assign io_d_unaligned = io_d_memrl == 2'h0 & _io_d_unaligned_T_10; // @[macros.scala 416:74]
endmodule
module muldiv(
  input         clock,
  input         reset,
  input         io_en,
  input  [4:0]  io_ctrl,
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_hi,
  output [31:0] io_lo,
  output        io_pending
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  _udiv_aclk; // @[muldiv.scala 193:23]
  wire  _udiv_s_axis_divisor_tvalid; // @[muldiv.scala 193:23]
  wire  _udiv_s_axis_divisor_tready; // @[muldiv.scala 193:23]
  wire [31:0] _udiv_s_axis_divisor_tdata; // @[muldiv.scala 193:23]
  wire  _udiv_s_axis_dividend_tvalid; // @[muldiv.scala 193:23]
  wire  _udiv_s_axis_dividend_tready; // @[muldiv.scala 193:23]
  wire [31:0] _udiv_s_axis_dividend_tdata; // @[muldiv.scala 193:23]
  wire  _udiv_m_axis_dout_tvalid; // @[muldiv.scala 193:23]
  wire [63:0] _udiv_m_axis_dout_tdata; // @[muldiv.scala 193:23]
  wire  _div_aclk; // @[muldiv.scala 205:23]
  wire  _div_s_axis_divisor_tvalid; // @[muldiv.scala 205:23]
  wire  _div_s_axis_divisor_tready; // @[muldiv.scala 205:23]
  wire [31:0] _div_s_axis_divisor_tdata; // @[muldiv.scala 205:23]
  wire  _div_s_axis_dividend_tvalid; // @[muldiv.scala 205:23]
  wire  _div_s_axis_dividend_tready; // @[muldiv.scala 205:23]
  wire [31:0] _div_s_axis_dividend_tdata; // @[muldiv.scala 205:23]
  wire  _div_m_axis_dout_tvalid; // @[muldiv.scala 205:23]
  wire [63:0] _div_m_axis_dout_tdata; // @[muldiv.scala 205:23]
  wire  _mul_CLK; // @[muldiv.scala 216:22]
  wire [31:0] _mul_A; // @[muldiv.scala 216:22]
  wire [31:0] _mul_B; // @[muldiv.scala 216:22]
  wire  _mul_CE; // @[muldiv.scala 216:22]
  wire [63:0] _mul_P; // @[muldiv.scala 216:22]
  wire  _umul_CLK; // @[muldiv.scala 226:23]
  wire [31:0] _umul_A; // @[muldiv.scala 226:23]
  wire [31:0] _umul_B; // @[muldiv.scala 226:23]
  wire  _umul_CE; // @[muldiv.scala 226:23]
  wire [63:0] _umul_P; // @[muldiv.scala 226:23]
  reg  counter_Reg; // @[muldiv.scala 82:30]
  reg  last_counter_Reg; // @[muldiv.scala 83:35]
  reg  in1_valid_u; // @[muldiv.scala 93:30]
  reg  in2_valid_u; // @[muldiv.scala 94:30]
  reg  in1_valid; // @[muldiv.scala 95:28]
  reg  in2_valid; // @[muldiv.scala 96:28]
  reg [31:0] a; // @[muldiv.scala 134:20]
  reg  b; // @[muldiv.scala 135:20]
  wire [5:0] _limit_T_1 = io_ctrl[0] ? 6'h22 : 6'h20; // @[muldiv.scala 137:17]
  wire [31:0] limit = {{26'd0}, _limit_T_1}; // @[muldiv.scala 136:21 137:11]
  wire [31:0] _a_T_3 = a + 32'h1; // @[muldiv.scala 138:55]
  reg [31:0] a_mul; // @[muldiv.scala 142:24]
  reg  b_mul; // @[muldiv.scala 143:24]
  wire  mul_counter_enable = io_en & (io_ctrl[2] | io_ctrl[3] | io_ctrl[4]); // @[muldiv.scala 145:43]
  wire [31:0] _a_mul_T_2 = 32'h3 - 32'h1; // @[muldiv.scala 148:68]
  wire  _a_mul_T_3 = a_mul == _a_mul_T_2; // @[muldiv.scala 148:54]
  wire [31:0] _a_mul_T_5 = a_mul + 32'h1; // @[muldiv.scala 148:85]
  wire  _T_2 = ~counter_Reg; // @[muldiv.scala 152:26]
  wire  in1_ready = _div_s_axis_dividend_tready; // @[muldiv.scala 103:24 212:15]
  wire  _GEN_0 = in1_ready | counter_Reg; // @[muldiv.scala 154:36 155:29 82:30]
  wire  in1_ready_u = _udiv_s_axis_dividend_tready; // @[muldiv.scala 101:26 200:17]
  wire  _GEN_1 = in1_ready_u | counter_Reg; // @[muldiv.scala 158:38 159:28 82:30]
  wire  _io_pending_T_8 = last_counter_Reg & _T_2 ? 1'h0 : 1'h1; // @[muldiv.scala 170:70]
  wire  _io_pending_T_16 = mul_counter_enable & b_mul; // @[muldiv.scala 171:12]
  wire [63:0] div_answer = _div_m_axis_dout_tdata; // @[muldiv.scala 118:27 213:16]
  wire [63:0] divu_answer = _udiv_m_axis_dout_tdata; // @[muldiv.scala 117:28 201:17]
  wire [63:0] mul_answer = _mul_P; // @[muldiv.scala 221:16 88:26]
  wire [63:0] mulu_answer = _umul_P; // @[muldiv.scala 231:17 87:27]
  wire [31:0] _io_lo_T_10 = io_ctrl[0] ? div_answer[63:32] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_lo_T_11 = io_ctrl[1] ? divu_answer[63:32] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_lo_T_12 = io_ctrl[2] ? mul_answer[31:0] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_lo_T_13 = io_ctrl[3] ? mulu_answer[31:0] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_lo_T_14 = io_ctrl[4] ? mulu_answer[31:0] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_lo_T_15 = _io_lo_T_10 | _io_lo_T_11; // @[Mux.scala 27:73]
  wire [31:0] _io_lo_T_16 = _io_lo_T_15 | _io_lo_T_12; // @[Mux.scala 27:73]
  wire [31:0] _io_lo_T_17 = _io_lo_T_16 | _io_lo_T_13; // @[Mux.scala 27:73]
  wire [31:0] _io_hi_T_10 = io_ctrl[0] ? div_answer[31:0] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_hi_T_11 = io_ctrl[1] ? divu_answer[31:0] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_hi_T_12 = io_ctrl[2] ? mul_answer[63:32] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_hi_T_13 = io_ctrl[3] ? mulu_answer[63:32] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_hi_T_14 = io_ctrl[4] ? mulu_answer[63:32] : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_hi_T_15 = _io_hi_T_10 | _io_hi_T_11; // @[Mux.scala 27:73]
  wire [31:0] _io_hi_T_16 = _io_hi_T_15 | _io_hi_T_12; // @[Mux.scala 27:73]
  wire [31:0] _io_hi_T_17 = _io_hi_T_16 | _io_hi_T_13; // @[Mux.scala 27:73]
  unsigned_div _udiv ( // @[muldiv.scala 193:23]
    .aclk(_udiv_aclk),
    .s_axis_divisor_tvalid(_udiv_s_axis_divisor_tvalid),
    .s_axis_divisor_tready(_udiv_s_axis_divisor_tready),
    .s_axis_divisor_tdata(_udiv_s_axis_divisor_tdata),
    .s_axis_dividend_tvalid(_udiv_s_axis_dividend_tvalid),
    .s_axis_dividend_tready(_udiv_s_axis_dividend_tready),
    .s_axis_dividend_tdata(_udiv_s_axis_dividend_tdata),
    .m_axis_dout_tvalid(_udiv_m_axis_dout_tvalid),
    .m_axis_dout_tdata(_udiv_m_axis_dout_tdata)
  );
  signed_div _div ( // @[muldiv.scala 205:23]
    .aclk(_div_aclk),
    .s_axis_divisor_tvalid(_div_s_axis_divisor_tvalid),
    .s_axis_divisor_tready(_div_s_axis_divisor_tready),
    .s_axis_divisor_tdata(_div_s_axis_divisor_tdata),
    .s_axis_dividend_tvalid(_div_s_axis_dividend_tvalid),
    .s_axis_dividend_tready(_div_s_axis_dividend_tready),
    .s_axis_dividend_tdata(_div_s_axis_dividend_tdata),
    .m_axis_dout_tvalid(_div_m_axis_dout_tvalid),
    .m_axis_dout_tdata(_div_m_axis_dout_tdata)
  );
  signed_mul _mul ( // @[muldiv.scala 216:22]
    .CLK(_mul_CLK),
    .A(_mul_A),
    .B(_mul_B),
    .CE(_mul_CE),
    .P(_mul_P)
  );
  unsigned_mul _umul ( // @[muldiv.scala 226:23]
    .CLK(_umul_CLK),
    .A(_umul_A),
    .B(_umul_B),
    .CE(_umul_CE),
    .P(_umul_P)
  );
  assign io_hi = _io_hi_T_17 | _io_hi_T_14; // @[Mux.scala 27:73]
  assign io_lo = _io_lo_T_17 | _io_lo_T_14; // @[Mux.scala 27:73]
  assign io_pending = io_en & (io_ctrl[0] | io_ctrl[1]) ? _io_pending_T_8 : _io_pending_T_16; // @[muldiv.scala 170:22]
  assign _udiv_aclk = clock; // @[muldiv.scala 194:19]
  assign _udiv_s_axis_divisor_tvalid = in2_valid_u; // @[muldiv.scala 195:36]
  assign _udiv_s_axis_divisor_tdata = io_en ? io_in2 : 32'h0; // @[muldiv.scala 112:23]
  assign _udiv_s_axis_dividend_tvalid = in1_valid_u; // @[muldiv.scala 197:37]
  assign _udiv_s_axis_dividend_tdata = io_en ? io_in1 : 32'h0; // @[muldiv.scala 113:24]
  assign _div_aclk = clock; // @[muldiv.scala 206:18]
  assign _div_s_axis_divisor_tvalid = in2_valid; // @[muldiv.scala 207:35]
  assign _div_s_axis_divisor_tdata = io_en ? io_in2 : 32'h0; // @[muldiv.scala 112:23]
  assign _div_s_axis_dividend_tvalid = in1_valid; // @[muldiv.scala 209:36]
  assign _div_s_axis_dividend_tdata = io_en ? io_in1 : 32'h0; // @[muldiv.scala 113:24]
  assign _mul_CLK = clock; // @[muldiv.scala 219:17]
  assign _mul_A = io_en ? io_in1 : 32'h0; // @[muldiv.scala 109:20]
  assign _mul_B = io_en ? io_in2 : 32'h0; // @[muldiv.scala 110:20]
  assign _mul_CE = io_en & (io_ctrl[2] | io_ctrl[3] | io_ctrl[4]); // @[muldiv.scala 145:43]
  assign _umul_CLK = clock; // @[muldiv.scala 229:18]
  assign _umul_A = io_en ? io_in1 : 32'h0; // @[muldiv.scala 109:20]
  assign _umul_B = io_en ? io_in2 : 32'h0; // @[muldiv.scala 110:20]
  assign _umul_CE = io_en & (io_ctrl[2] | io_ctrl[3] | io_ctrl[4]); // @[muldiv.scala 145:43]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[muldiv.scala 152:47]
      counter_Reg <= 1'h0; // @[muldiv.scala 153:27 157:31 82:30]
    end else if (io_en & ~counter_Reg) begin // @[muldiv.scala 163:24]
      if (io_ctrl[0]) begin // @[muldiv.scala 165:25]
        counter_Reg <= _GEN_0;
      end else if (io_ctrl[1]) begin
        counter_Reg <= _GEN_1;
      end
    end else if (b) begin // @[muldiv.scala 82:30]
      counter_Reg <= 1'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[muldiv.scala 83:35]
      last_counter_Reg <= 1'h0; // @[muldiv.scala 83:35]
    end else begin
      last_counter_Reg <= counter_Reg; // @[muldiv.scala 84:22]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[muldiv.scala 93:30]
      in1_valid_u <= 1'h0; // @[muldiv.scala 93:30]
    end else begin
      in1_valid_u <= 1'h1; // @[muldiv.scala 122:17]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[muldiv.scala 94:30]
      in2_valid_u <= 1'h0; // @[muldiv.scala 94:30]
    end else begin
      in2_valid_u <= 1'h1; // @[muldiv.scala 123:17]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[muldiv.scala 95:28]
      in1_valid <= 1'h0; // @[muldiv.scala 95:28]
    end else begin
      in1_valid <= 1'h1; // @[muldiv.scala 120:15]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[muldiv.scala 96:28]
      in2_valid <= 1'h0; // @[muldiv.scala 96:28]
    end else begin
      in2_valid <= 1'h1; // @[muldiv.scala 121:15]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[muldiv.scala 138:13]
      a <= 32'h0; // @[muldiv.scala 138:36]
    end else if (counter_Reg) begin
      if (a == limit) begin
        a <= 32'h0;
      end else begin
        a <= _a_T_3;
      end
    end else begin
      a <= 32'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[muldiv.scala 139:16]
      b <= 1'h0;
    end else begin
      b <= a == limit;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[muldiv.scala 148:17]
      a_mul <= 32'h0; // @[muldiv.scala 148:47]
    end else if (mul_counter_enable) begin
      if (a_mul == _a_mul_T_2) begin
        a_mul <= 32'h0;
      end else begin
        a_mul <= _a_mul_T_5;
      end
    end else begin
      a_mul <= 32'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[muldiv.scala 149:17]
      b_mul <= 1'h0;
    end else if (_a_mul_T_3) begin
      b_mul <= 1'h0;
    end else begin
      b_mul <= 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counter_Reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  last_counter_Reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in1_valid_u = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in2_valid_u = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  in1_valid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  in2_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  a = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  b = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  a_mul = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  b_mul = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    counter_Reg = 1'h0;
  end
  if (reset) begin
    last_counter_Reg = 1'h0;
  end
  if (reset) begin
    in1_valid_u = 1'h0;
  end
  if (reset) begin
    in2_valid_u = 1'h0;
  end
  if (reset) begin
    in1_valid = 1'h0;
  end
  if (reset) begin
    in2_valid = 1'h0;
  end
  if (reset) begin
    a = 32'h0;
  end
  if (reset) begin
    b = 1'h0;
  end
  if (reset) begin
    a_mul = 32'h0;
  end
  if (reset) begin
    b_mul = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module regfile(
  input         clock,
  input         reset,
  input  [4:0]  io_A1,
  input  [4:0]  io_A2,
  input         io_WE3,
  input  [4:0]  io_A3,
  input  [31:0] io_WD3,
  output [31:0] io_RD1,
  output [31:0] io_RD2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0; // @[regfile.scala 23:23]
  reg [31:0] regs_1; // @[regfile.scala 23:23]
  reg [31:0] regs_2; // @[regfile.scala 23:23]
  reg [31:0] regs_3; // @[regfile.scala 23:23]
  reg [31:0] regs_4; // @[regfile.scala 23:23]
  reg [31:0] regs_5; // @[regfile.scala 23:23]
  reg [31:0] regs_6; // @[regfile.scala 23:23]
  reg [31:0] regs_7; // @[regfile.scala 23:23]
  reg [31:0] regs_8; // @[regfile.scala 23:23]
  reg [31:0] regs_9; // @[regfile.scala 23:23]
  reg [31:0] regs_10; // @[regfile.scala 23:23]
  reg [31:0] regs_11; // @[regfile.scala 23:23]
  reg [31:0] regs_12; // @[regfile.scala 23:23]
  reg [31:0] regs_13; // @[regfile.scala 23:23]
  reg [31:0] regs_14; // @[regfile.scala 23:23]
  reg [31:0] regs_15; // @[regfile.scala 23:23]
  reg [31:0] regs_16; // @[regfile.scala 23:23]
  reg [31:0] regs_17; // @[regfile.scala 23:23]
  reg [31:0] regs_18; // @[regfile.scala 23:23]
  reg [31:0] regs_19; // @[regfile.scala 23:23]
  reg [31:0] regs_20; // @[regfile.scala 23:23]
  reg [31:0] regs_21; // @[regfile.scala 23:23]
  reg [31:0] regs_22; // @[regfile.scala 23:23]
  reg [31:0] regs_23; // @[regfile.scala 23:23]
  reg [31:0] regs_24; // @[regfile.scala 23:23]
  reg [31:0] regs_25; // @[regfile.scala 23:23]
  reg [31:0] regs_26; // @[regfile.scala 23:23]
  reg [31:0] regs_27; // @[regfile.scala 23:23]
  reg [31:0] regs_28; // @[regfile.scala 23:23]
  reg [31:0] regs_29; // @[regfile.scala 23:23]
  reg [31:0] regs_30; // @[regfile.scala 23:23]
  reg [31:0] regs_31; // @[regfile.scala 23:23]
  wire [31:0] _GEN_1 = 5'h1 == io_A3 ? regs_1 : regs_0; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_2 = 5'h2 == io_A3 ? regs_2 : _GEN_1; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_3 = 5'h3 == io_A3 ? regs_3 : _GEN_2; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_4 = 5'h4 == io_A3 ? regs_4 : _GEN_3; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_5 = 5'h5 == io_A3 ? regs_5 : _GEN_4; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_6 = 5'h6 == io_A3 ? regs_6 : _GEN_5; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_7 = 5'h7 == io_A3 ? regs_7 : _GEN_6; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_8 = 5'h8 == io_A3 ? regs_8 : _GEN_7; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_9 = 5'h9 == io_A3 ? regs_9 : _GEN_8; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_10 = 5'ha == io_A3 ? regs_10 : _GEN_9; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_11 = 5'hb == io_A3 ? regs_11 : _GEN_10; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_12 = 5'hc == io_A3 ? regs_12 : _GEN_11; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_13 = 5'hd == io_A3 ? regs_13 : _GEN_12; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_14 = 5'he == io_A3 ? regs_14 : _GEN_13; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_15 = 5'hf == io_A3 ? regs_15 : _GEN_14; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_16 = 5'h10 == io_A3 ? regs_16 : _GEN_15; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_17 = 5'h11 == io_A3 ? regs_17 : _GEN_16; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_18 = 5'h12 == io_A3 ? regs_18 : _GEN_17; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_19 = 5'h13 == io_A3 ? regs_19 : _GEN_18; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_20 = 5'h14 == io_A3 ? regs_20 : _GEN_19; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_21 = 5'h15 == io_A3 ? regs_21 : _GEN_20; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_22 = 5'h16 == io_A3 ? regs_22 : _GEN_21; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_23 = 5'h17 == io_A3 ? regs_23 : _GEN_22; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_24 = 5'h18 == io_A3 ? regs_24 : _GEN_23; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_25 = 5'h19 == io_A3 ? regs_25 : _GEN_24; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_26 = 5'h1a == io_A3 ? regs_26 : _GEN_25; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_27 = 5'h1b == io_A3 ? regs_27 : _GEN_26; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_28 = 5'h1c == io_A3 ? regs_28 : _GEN_27; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_29 = 5'h1d == io_A3 ? regs_29 : _GEN_28; // @[regfile.scala 25:{23,23}]
  wire [31:0] _GEN_65 = 5'h1 == io_A1 ? regs_1 : regs_0; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_66 = 5'h2 == io_A1 ? regs_2 : _GEN_65; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_67 = 5'h3 == io_A1 ? regs_3 : _GEN_66; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_68 = 5'h4 == io_A1 ? regs_4 : _GEN_67; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_69 = 5'h5 == io_A1 ? regs_5 : _GEN_68; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_70 = 5'h6 == io_A1 ? regs_6 : _GEN_69; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_71 = 5'h7 == io_A1 ? regs_7 : _GEN_70; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_72 = 5'h8 == io_A1 ? regs_8 : _GEN_71; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_73 = 5'h9 == io_A1 ? regs_9 : _GEN_72; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_74 = 5'ha == io_A1 ? regs_10 : _GEN_73; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_75 = 5'hb == io_A1 ? regs_11 : _GEN_74; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_76 = 5'hc == io_A1 ? regs_12 : _GEN_75; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_77 = 5'hd == io_A1 ? regs_13 : _GEN_76; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_78 = 5'he == io_A1 ? regs_14 : _GEN_77; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_79 = 5'hf == io_A1 ? regs_15 : _GEN_78; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_80 = 5'h10 == io_A1 ? regs_16 : _GEN_79; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_81 = 5'h11 == io_A1 ? regs_17 : _GEN_80; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_82 = 5'h12 == io_A1 ? regs_18 : _GEN_81; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_83 = 5'h13 == io_A1 ? regs_19 : _GEN_82; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_84 = 5'h14 == io_A1 ? regs_20 : _GEN_83; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_85 = 5'h15 == io_A1 ? regs_21 : _GEN_84; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_86 = 5'h16 == io_A1 ? regs_22 : _GEN_85; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_87 = 5'h17 == io_A1 ? regs_23 : _GEN_86; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_88 = 5'h18 == io_A1 ? regs_24 : _GEN_87; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_89 = 5'h19 == io_A1 ? regs_25 : _GEN_88; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_90 = 5'h1a == io_A1 ? regs_26 : _GEN_89; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_91 = 5'h1b == io_A1 ? regs_27 : _GEN_90; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_92 = 5'h1c == io_A1 ? regs_28 : _GEN_91; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_93 = 5'h1d == io_A1 ? regs_29 : _GEN_92; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_94 = 5'h1e == io_A1 ? regs_30 : _GEN_93; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_95 = 5'h1f == io_A1 ? regs_31 : _GEN_94; // @[regfile.scala 34:{19,19}]
  wire [31:0] _GEN_97 = 5'h1 == io_A2 ? regs_1 : regs_0; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_98 = 5'h2 == io_A2 ? regs_2 : _GEN_97; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_99 = 5'h3 == io_A2 ? regs_3 : _GEN_98; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_100 = 5'h4 == io_A2 ? regs_4 : _GEN_99; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_101 = 5'h5 == io_A2 ? regs_5 : _GEN_100; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_102 = 5'h6 == io_A2 ? regs_6 : _GEN_101; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_103 = 5'h7 == io_A2 ? regs_7 : _GEN_102; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_104 = 5'h8 == io_A2 ? regs_8 : _GEN_103; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_105 = 5'h9 == io_A2 ? regs_9 : _GEN_104; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_106 = 5'ha == io_A2 ? regs_10 : _GEN_105; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_107 = 5'hb == io_A2 ? regs_11 : _GEN_106; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_108 = 5'hc == io_A2 ? regs_12 : _GEN_107; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_109 = 5'hd == io_A2 ? regs_13 : _GEN_108; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_110 = 5'he == io_A2 ? regs_14 : _GEN_109; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_111 = 5'hf == io_A2 ? regs_15 : _GEN_110; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_112 = 5'h10 == io_A2 ? regs_16 : _GEN_111; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_113 = 5'h11 == io_A2 ? regs_17 : _GEN_112; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_114 = 5'h12 == io_A2 ? regs_18 : _GEN_113; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_115 = 5'h13 == io_A2 ? regs_19 : _GEN_114; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_116 = 5'h14 == io_A2 ? regs_20 : _GEN_115; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_117 = 5'h15 == io_A2 ? regs_21 : _GEN_116; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_118 = 5'h16 == io_A2 ? regs_22 : _GEN_117; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_119 = 5'h17 == io_A2 ? regs_23 : _GEN_118; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_120 = 5'h18 == io_A2 ? regs_24 : _GEN_119; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_121 = 5'h19 == io_A2 ? regs_25 : _GEN_120; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_122 = 5'h1a == io_A2 ? regs_26 : _GEN_121; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_123 = 5'h1b == io_A2 ? regs_27 : _GEN_122; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_124 = 5'h1c == io_A2 ? regs_28 : _GEN_123; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_125 = 5'h1d == io_A2 ? regs_29 : _GEN_124; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_126 = 5'h1e == io_A2 ? regs_30 : _GEN_125; // @[regfile.scala 35:{19,19}]
  wire [31:0] _GEN_127 = 5'h1f == io_A2 ? regs_31 : _GEN_126; // @[regfile.scala 35:{19,19}]
  assign io_RD1 = io_WE3 & io_A1 == io_A3 ? io_WD3 : _GEN_95; // @[regfile.scala 34:19]
  assign io_RD2 = io_WE3 & io_A2 == io_A3 ? io_WD3 : _GEN_127; // @[regfile.scala 35:19]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_0 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h0 == io_A3) begin // @[regfile.scala 24:13]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_0 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_0 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_0 <= regs_30;
      end else begin
        regs_0 <= _GEN_29;
      end
    end else begin
      regs_0 <= 32'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_1 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h1 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_1 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_1 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_1 <= regs_30;
      end else begin
        regs_1 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_2 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h2 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_2 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_2 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_2 <= regs_30;
      end else begin
        regs_2 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_3 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h3 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_3 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_3 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_3 <= regs_30;
      end else begin
        regs_3 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_4 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h4 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_4 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_4 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_4 <= regs_30;
      end else begin
        regs_4 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_5 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h5 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_5 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_5 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_5 <= regs_30;
      end else begin
        regs_5 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_6 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h6 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_6 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_6 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_6 <= regs_30;
      end else begin
        regs_6 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_7 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h7 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_7 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_7 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_7 <= regs_30;
      end else begin
        regs_7 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_8 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h8 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_8 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_8 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_8 <= regs_30;
      end else begin
        regs_8 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_9 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h9 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_9 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_9 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_9 <= regs_30;
      end else begin
        regs_9 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_10 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'ha == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_10 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_10 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_10 <= regs_30;
      end else begin
        regs_10 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_11 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'hb == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_11 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_11 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_11 <= regs_30;
      end else begin
        regs_11 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_12 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'hc == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_12 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_12 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_12 <= regs_30;
      end else begin
        regs_12 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_13 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'hd == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_13 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_13 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_13 <= regs_30;
      end else begin
        regs_13 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_14 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'he == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_14 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_14 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_14 <= regs_30;
      end else begin
        regs_14 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_15 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'hf == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_15 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_15 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_15 <= regs_30;
      end else begin
        regs_15 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_16 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h10 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_16 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_16 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_16 <= regs_30;
      end else begin
        regs_16 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_17 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h11 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_17 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_17 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_17 <= regs_30;
      end else begin
        regs_17 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_18 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h12 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_18 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_18 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_18 <= regs_30;
      end else begin
        regs_18 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_19 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h13 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_19 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_19 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_19 <= regs_30;
      end else begin
        regs_19 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_20 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h14 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_20 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_20 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_20 <= regs_30;
      end else begin
        regs_20 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_21 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h15 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_21 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_21 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_21 <= regs_30;
      end else begin
        regs_21 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_22 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h16 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_22 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_22 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_22 <= regs_30;
      end else begin
        regs_22 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_23 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h17 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_23 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_23 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_23 <= regs_30;
      end else begin
        regs_23 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_24 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h18 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_24 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_24 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_24 <= regs_30;
      end else begin
        regs_24 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_25 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h19 == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_25 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_25 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_25 <= regs_30;
      end else begin
        regs_25 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_26 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h1a == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_26 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_26 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_26 <= regs_30;
      end else begin
        regs_26 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_27 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h1b == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_27 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_27 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_27 <= regs_30;
      end else begin
        regs_27 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_28 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h1c == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_28 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_28 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_28 <= regs_30;
      end else begin
        regs_28 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_29 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h1d == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_29 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_29 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_29 <= regs_30;
      end else begin
        regs_29 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_30 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h1e == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_30 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_30 <= regs_31;
      end else if (!(5'h1e == io_A3)) begin
        regs_30 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 25:17]
      regs_31 <= 32'h0; // @[regfile.scala 25:{23,23,23,23,23}]
    end else if (5'h1f == io_A3) begin // @[regfile.scala 23:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_31 <= io_WD3;
      end else if (!(5'h1f == io_A3)) begin
        if (5'h1e == io_A3) begin
          regs_31 <= regs_30;
        end else begin
          regs_31 <= _GEN_29;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    regs_0 = 32'h0;
  end
  if (reset) begin
    regs_1 = 32'h0;
  end
  if (reset) begin
    regs_2 = 32'h0;
  end
  if (reset) begin
    regs_3 = 32'h0;
  end
  if (reset) begin
    regs_4 = 32'h0;
  end
  if (reset) begin
    regs_5 = 32'h0;
  end
  if (reset) begin
    regs_6 = 32'h0;
  end
  if (reset) begin
    regs_7 = 32'h0;
  end
  if (reset) begin
    regs_8 = 32'h0;
  end
  if (reset) begin
    regs_9 = 32'h0;
  end
  if (reset) begin
    regs_10 = 32'h0;
  end
  if (reset) begin
    regs_11 = 32'h0;
  end
  if (reset) begin
    regs_12 = 32'h0;
  end
  if (reset) begin
    regs_13 = 32'h0;
  end
  if (reset) begin
    regs_14 = 32'h0;
  end
  if (reset) begin
    regs_15 = 32'h0;
  end
  if (reset) begin
    regs_16 = 32'h0;
  end
  if (reset) begin
    regs_17 = 32'h0;
  end
  if (reset) begin
    regs_18 = 32'h0;
  end
  if (reset) begin
    regs_19 = 32'h0;
  end
  if (reset) begin
    regs_20 = 32'h0;
  end
  if (reset) begin
    regs_21 = 32'h0;
  end
  if (reset) begin
    regs_22 = 32'h0;
  end
  if (reset) begin
    regs_23 = 32'h0;
  end
  if (reset) begin
    regs_24 = 32'h0;
  end
  if (reset) begin
    regs_25 = 32'h0;
  end
  if (reset) begin
    regs_26 = 32'h0;
  end
  if (reset) begin
    regs_27 = 32'h0;
  end
  if (reset) begin
    regs_28 = 32'h0;
  end
  if (reset) begin
    regs_29 = 32'h0;
  end
  if (reset) begin
    regs_30 = 32'h0;
  end
  if (reset) begin
    regs_31 = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Look_up_table_read_first_(
  input          clock,
  input          reset,
  input  [3:0]   io_ar_addr,
  input  [3:0]   io_aw_addr,
  input          io_write,
  input  [135:0] io_in,
  output [135:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [159:0] _RAND_4;
  reg [159:0] _RAND_5;
  reg [159:0] _RAND_6;
  reg [159:0] _RAND_7;
  reg [159:0] _RAND_8;
  reg [159:0] _RAND_9;
  reg [159:0] _RAND_10;
  reg [159:0] _RAND_11;
  reg [159:0] _RAND_12;
  reg [159:0] _RAND_13;
  reg [159:0] _RAND_14;
  reg [159:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [135:0] btb_0; // @[ports_lookup_table.scala 81:22]
  reg [135:0] btb_1; // @[ports_lookup_table.scala 81:22]
  reg [135:0] btb_2; // @[ports_lookup_table.scala 81:22]
  reg [135:0] btb_3; // @[ports_lookup_table.scala 81:22]
  reg [135:0] btb_4; // @[ports_lookup_table.scala 81:22]
  reg [135:0] btb_5; // @[ports_lookup_table.scala 81:22]
  reg [135:0] btb_6; // @[ports_lookup_table.scala 81:22]
  reg [135:0] btb_7; // @[ports_lookup_table.scala 81:22]
  reg [135:0] btb_8; // @[ports_lookup_table.scala 81:22]
  reg [135:0] btb_9; // @[ports_lookup_table.scala 81:22]
  reg [135:0] btb_10; // @[ports_lookup_table.scala 81:22]
  reg [135:0] btb_11; // @[ports_lookup_table.scala 81:22]
  reg [135:0] btb_12; // @[ports_lookup_table.scala 81:22]
  reg [135:0] btb_13; // @[ports_lookup_table.scala 81:22]
  reg [135:0] btb_14; // @[ports_lookup_table.scala 81:22]
  reg [135:0] btb_15; // @[ports_lookup_table.scala 81:22]
  wire [135:0] _GEN_1 = 4'h1 == io_ar_addr ? btb_1 : btb_0; // @[ports_lookup_table.scala 82:{12,12}]
  wire [135:0] _GEN_2 = 4'h2 == io_ar_addr ? btb_2 : _GEN_1; // @[ports_lookup_table.scala 82:{12,12}]
  wire [135:0] _GEN_3 = 4'h3 == io_ar_addr ? btb_3 : _GEN_2; // @[ports_lookup_table.scala 82:{12,12}]
  wire [135:0] _GEN_4 = 4'h4 == io_ar_addr ? btb_4 : _GEN_3; // @[ports_lookup_table.scala 82:{12,12}]
  wire [135:0] _GEN_5 = 4'h5 == io_ar_addr ? btb_5 : _GEN_4; // @[ports_lookup_table.scala 82:{12,12}]
  wire [135:0] _GEN_6 = 4'h6 == io_ar_addr ? btb_6 : _GEN_5; // @[ports_lookup_table.scala 82:{12,12}]
  wire [135:0] _GEN_7 = 4'h7 == io_ar_addr ? btb_7 : _GEN_6; // @[ports_lookup_table.scala 82:{12,12}]
  wire [135:0] _GEN_8 = 4'h8 == io_ar_addr ? btb_8 : _GEN_7; // @[ports_lookup_table.scala 82:{12,12}]
  wire [135:0] _GEN_9 = 4'h9 == io_ar_addr ? btb_9 : _GEN_8; // @[ports_lookup_table.scala 82:{12,12}]
  wire [135:0] _GEN_10 = 4'ha == io_ar_addr ? btb_10 : _GEN_9; // @[ports_lookup_table.scala 82:{12,12}]
  wire [135:0] _GEN_11 = 4'hb == io_ar_addr ? btb_11 : _GEN_10; // @[ports_lookup_table.scala 82:{12,12}]
  wire [135:0] _GEN_12 = 4'hc == io_ar_addr ? btb_12 : _GEN_11; // @[ports_lookup_table.scala 82:{12,12}]
  wire [135:0] _GEN_13 = 4'hd == io_ar_addr ? btb_13 : _GEN_12; // @[ports_lookup_table.scala 82:{12,12}]
  wire [135:0] _GEN_14 = 4'he == io_ar_addr ? btb_14 : _GEN_13; // @[ports_lookup_table.scala 82:{12,12}]
  wire [135:0] _GEN_17 = 4'h1 == io_aw_addr ? btb_1 : btb_0; // @[ports_lookup_table.scala 83:{27,27}]
  wire [135:0] _GEN_18 = 4'h2 == io_aw_addr ? btb_2 : _GEN_17; // @[ports_lookup_table.scala 83:{27,27}]
  wire [135:0] _GEN_19 = 4'h3 == io_aw_addr ? btb_3 : _GEN_18; // @[ports_lookup_table.scala 83:{27,27}]
  wire [135:0] _GEN_20 = 4'h4 == io_aw_addr ? btb_4 : _GEN_19; // @[ports_lookup_table.scala 83:{27,27}]
  wire [135:0] _GEN_21 = 4'h5 == io_aw_addr ? btb_5 : _GEN_20; // @[ports_lookup_table.scala 83:{27,27}]
  wire [135:0] _GEN_22 = 4'h6 == io_aw_addr ? btb_6 : _GEN_21; // @[ports_lookup_table.scala 83:{27,27}]
  wire [135:0] _GEN_23 = 4'h7 == io_aw_addr ? btb_7 : _GEN_22; // @[ports_lookup_table.scala 83:{27,27}]
  wire [135:0] _GEN_24 = 4'h8 == io_aw_addr ? btb_8 : _GEN_23; // @[ports_lookup_table.scala 83:{27,27}]
  wire [135:0] _GEN_25 = 4'h9 == io_aw_addr ? btb_9 : _GEN_24; // @[ports_lookup_table.scala 83:{27,27}]
  wire [135:0] _GEN_26 = 4'ha == io_aw_addr ? btb_10 : _GEN_25; // @[ports_lookup_table.scala 83:{27,27}]
  wire [135:0] _GEN_27 = 4'hb == io_aw_addr ? btb_11 : _GEN_26; // @[ports_lookup_table.scala 83:{27,27}]
  wire [135:0] _GEN_28 = 4'hc == io_aw_addr ? btb_12 : _GEN_27; // @[ports_lookup_table.scala 83:{27,27}]
  wire [135:0] _GEN_29 = 4'hd == io_aw_addr ? btb_13 : _GEN_28; // @[ports_lookup_table.scala 83:{27,27}]
  assign io_out = 4'hf == io_ar_addr ? btb_15 : _GEN_14; // @[ports_lookup_table.scala 82:{12,12}]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_0 <= 136'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_0 <= io_in;
      end else if (4'hf == io_aw_addr) begin
        btb_0 <= btb_15;
      end else if (4'he == io_aw_addr) begin
        btb_0 <= btb_14;
      end else begin
        btb_0 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_1 <= 136'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_1 <= io_in;
      end else if (4'hf == io_aw_addr) begin
        btb_1 <= btb_15;
      end else if (4'he == io_aw_addr) begin
        btb_1 <= btb_14;
      end else begin
        btb_1 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_2 <= 136'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_2 <= io_in;
      end else if (4'hf == io_aw_addr) begin
        btb_2 <= btb_15;
      end else if (4'he == io_aw_addr) begin
        btb_2 <= btb_14;
      end else begin
        btb_2 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_3 <= 136'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_3 <= io_in;
      end else if (4'hf == io_aw_addr) begin
        btb_3 <= btb_15;
      end else if (4'he == io_aw_addr) begin
        btb_3 <= btb_14;
      end else begin
        btb_3 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_4 <= 136'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_4 <= io_in;
      end else if (4'hf == io_aw_addr) begin
        btb_4 <= btb_15;
      end else if (4'he == io_aw_addr) begin
        btb_4 <= btb_14;
      end else begin
        btb_4 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_5 <= 136'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_5 <= io_in;
      end else if (4'hf == io_aw_addr) begin
        btb_5 <= btb_15;
      end else if (4'he == io_aw_addr) begin
        btb_5 <= btb_14;
      end else begin
        btb_5 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_6 <= 136'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_6 <= io_in;
      end else if (4'hf == io_aw_addr) begin
        btb_6 <= btb_15;
      end else if (4'he == io_aw_addr) begin
        btb_6 <= btb_14;
      end else begin
        btb_6 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_7 <= 136'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_7 <= io_in;
      end else if (4'hf == io_aw_addr) begin
        btb_7 <= btb_15;
      end else if (4'he == io_aw_addr) begin
        btb_7 <= btb_14;
      end else begin
        btb_7 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_8 <= 136'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_8 <= io_in;
      end else if (4'hf == io_aw_addr) begin
        btb_8 <= btb_15;
      end else if (4'he == io_aw_addr) begin
        btb_8 <= btb_14;
      end else begin
        btb_8 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_9 <= 136'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_9 <= io_in;
      end else if (4'hf == io_aw_addr) begin
        btb_9 <= btb_15;
      end else if (4'he == io_aw_addr) begin
        btb_9 <= btb_14;
      end else begin
        btb_9 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_10 <= 136'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_10 <= io_in;
      end else if (4'hf == io_aw_addr) begin
        btb_10 <= btb_15;
      end else if (4'he == io_aw_addr) begin
        btb_10 <= btb_14;
      end else begin
        btb_10 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_11 <= 136'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_11 <= io_in;
      end else if (4'hf == io_aw_addr) begin
        btb_11 <= btb_15;
      end else if (4'he == io_aw_addr) begin
        btb_11 <= btb_14;
      end else begin
        btb_11 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_12 <= 136'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_12 <= io_in;
      end else if (4'hf == io_aw_addr) begin
        btb_12 <= btb_15;
      end else if (4'he == io_aw_addr) begin
        btb_12 <= btb_14;
      end else begin
        btb_12 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_13 <= 136'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_13 <= io_in;
      end else if (4'hf == io_aw_addr) begin
        btb_13 <= btb_15;
      end else if (4'he == io_aw_addr) begin
        btb_13 <= btb_14;
      end else begin
        btb_13 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_14 <= 136'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_14 <= io_in;
      end else if (4'hf == io_aw_addr) begin
        btb_14 <= btb_15;
      end else if (!(4'he == io_aw_addr)) begin
        btb_14 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_15 <= 136'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_15 <= io_in;
      end else if (!(4'hf == io_aw_addr)) begin
        if (4'he == io_aw_addr) begin
          btb_15 <= btb_14;
        end else begin
          btb_15 <= _GEN_29;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{`RANDOM}};
  btb_0 = _RAND_0[135:0];
  _RAND_1 = {5{`RANDOM}};
  btb_1 = _RAND_1[135:0];
  _RAND_2 = {5{`RANDOM}};
  btb_2 = _RAND_2[135:0];
  _RAND_3 = {5{`RANDOM}};
  btb_3 = _RAND_3[135:0];
  _RAND_4 = {5{`RANDOM}};
  btb_4 = _RAND_4[135:0];
  _RAND_5 = {5{`RANDOM}};
  btb_5 = _RAND_5[135:0];
  _RAND_6 = {5{`RANDOM}};
  btb_6 = _RAND_6[135:0];
  _RAND_7 = {5{`RANDOM}};
  btb_7 = _RAND_7[135:0];
  _RAND_8 = {5{`RANDOM}};
  btb_8 = _RAND_8[135:0];
  _RAND_9 = {5{`RANDOM}};
  btb_9 = _RAND_9[135:0];
  _RAND_10 = {5{`RANDOM}};
  btb_10 = _RAND_10[135:0];
  _RAND_11 = {5{`RANDOM}};
  btb_11 = _RAND_11[135:0];
  _RAND_12 = {5{`RANDOM}};
  btb_12 = _RAND_12[135:0];
  _RAND_13 = {5{`RANDOM}};
  btb_13 = _RAND_13[135:0];
  _RAND_14 = {5{`RANDOM}};
  btb_14 = _RAND_14[135:0];
  _RAND_15 = {5{`RANDOM}};
  btb_15 = _RAND_15[135:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    btb_0 = 136'h0;
  end
  if (reset) begin
    btb_1 = 136'h0;
  end
  if (reset) begin
    btb_2 = 136'h0;
  end
  if (reset) begin
    btb_3 = 136'h0;
  end
  if (reset) begin
    btb_4 = 136'h0;
  end
  if (reset) begin
    btb_5 = 136'h0;
  end
  if (reset) begin
    btb_6 = 136'h0;
  end
  if (reset) begin
    btb_7 = 136'h0;
  end
  if (reset) begin
    btb_8 = 136'h0;
  end
  if (reset) begin
    btb_9 = 136'h0;
  end
  if (reset) begin
    btb_10 = 136'h0;
  end
  if (reset) begin
    btb_11 = 136'h0;
  end
  if (reset) begin
    btb_12 = 136'h0;
  end
  if (reset) begin
    btb_13 = 136'h0;
  end
  if (reset) begin
    btb_14 = 136'h0;
  end
  if (reset) begin
    btb_15 = 136'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module fifo(
  input          clock,
  input          reset,
  input  [1:0]   io_read_en,
  input  [1:0]   io_write_en,
  output [135:0] io_read_out_0,
  input  [135:0] io_write_in_0,
  output         io_full,
  output         io_empty,
  input          io_point_write_en,
  input          io_point_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  Look_up_table_read_first__clock; // @[fifo.scala 42:55]
  wire  Look_up_table_read_first__reset; // @[fifo.scala 42:55]
  wire [3:0] Look_up_table_read_first__io_ar_addr; // @[fifo.scala 42:55]
  wire [3:0] Look_up_table_read_first__io_aw_addr; // @[fifo.scala 42:55]
  wire  Look_up_table_read_first__io_write; // @[fifo.scala 42:55]
  wire [135:0] Look_up_table_read_first__io_in; // @[fifo.scala 42:55]
  wire [135:0] Look_up_table_read_first__io_out; // @[fifo.scala 42:55]
  wire  Look_up_table_read_first__1_clock; // @[fifo.scala 42:55]
  wire  Look_up_table_read_first__1_reset; // @[fifo.scala 42:55]
  wire [3:0] Look_up_table_read_first__1_io_ar_addr; // @[fifo.scala 42:55]
  wire [3:0] Look_up_table_read_first__1_io_aw_addr; // @[fifo.scala 42:55]
  wire  Look_up_table_read_first__1_io_write; // @[fifo.scala 42:55]
  wire [135:0] Look_up_table_read_first__1_io_in; // @[fifo.scala 42:55]
  wire [135:0] Look_up_table_read_first__1_io_out; // @[fifo.scala 42:55]
  wire  Look_up_table_read_first__2_clock; // @[fifo.scala 42:55]
  wire  Look_up_table_read_first__2_reset; // @[fifo.scala 42:55]
  wire [3:0] Look_up_table_read_first__2_io_ar_addr; // @[fifo.scala 42:55]
  wire [3:0] Look_up_table_read_first__2_io_aw_addr; // @[fifo.scala 42:55]
  wire  Look_up_table_read_first__2_io_write; // @[fifo.scala 42:55]
  wire [135:0] Look_up_table_read_first__2_io_in; // @[fifo.scala 42:55]
  wire [135:0] Look_up_table_read_first__2_io_out; // @[fifo.scala 42:55]
  wire  Look_up_table_read_first__3_clock; // @[fifo.scala 42:55]
  wire  Look_up_table_read_first__3_reset; // @[fifo.scala 42:55]
  wire [3:0] Look_up_table_read_first__3_io_ar_addr; // @[fifo.scala 42:55]
  wire [3:0] Look_up_table_read_first__3_io_aw_addr; // @[fifo.scala 42:55]
  wire  Look_up_table_read_first__3_io_write; // @[fifo.scala 42:55]
  wire [135:0] Look_up_table_read_first__3_io_in; // @[fifo.scala 42:55]
  wire [135:0] Look_up_table_read_first__3_io_out; // @[fifo.scala 42:55]
  reg [1:0] write_banks_points; // @[fifo.scala 43:37]
  reg [3:0] write_length_points; // @[fifo.scala 44:38]
  reg [1:0] read_banks_points; // @[fifo.scala 45:36]
  reg [3:0] read_length_points; // @[fifo.scala 46:37]
  wire  _fifo_banks_3_write_T_1 = write_banks_points == 2'h3; // @[Mux.scala 81:61]
  wire  point_write_tag = io_point_write_en & (~io_empty | io_empty & io_write_en != 2'h0); // @[fifo.scala 87:49]
  wire [1:0] _write_banks_points_T_2 = read_banks_points + 2'h1; // @[fifo.scala 93:95]
  wire [1:0] _write_banks_points_T_4 = write_banks_points + io_write_en; // @[fifo.scala 93:121]
  wire [3:0] _GEN_4 = {{3'd0}, read_banks_points == 2'h3}; // @[fifo.scala 97:97]
  wire [3:0] _write_length_points_T_4 = read_length_points + _GEN_4; // @[fifo.scala 97:97]
  wire [2:0] _write_length_points_T_5 = {1'h0,write_banks_points}; // @[Cat.scala 31:58]
  wire [2:0] _GEN_5 = {{1'd0}, io_write_en}; // @[fifo.scala 97:200]
  wire [2:0] _write_length_points_T_7 = _write_length_points_T_5 + _GEN_5; // @[fifo.scala 97:200]
  wire [3:0] _GEN_6 = {{3'd0}, _write_length_points_T_7[2]}; // @[fifo.scala 97:159]
  wire [3:0] _write_length_points_T_11 = write_length_points + _GEN_6; // @[fifo.scala 97:159]
  wire [1:0] _read_banks_points_T_1 = read_banks_points + io_read_en; // @[fifo.scala 98:68]
  wire [2:0] _read_length_points_T = {1'h0,read_banks_points}; // @[Cat.scala 31:58]
  wire [2:0] _GEN_7 = {{1'd0}, io_read_en}; // @[fifo.scala 99:110]
  wire [2:0] _read_length_points_T_2 = _read_length_points_T + _GEN_7; // @[fifo.scala 99:110]
  wire [3:0] _GEN_8 = {{3'd0}, _read_length_points_T_2[2]}; // @[fifo.scala 99:71]
  wire [3:0] _read_length_points_T_6 = read_length_points + _GEN_8; // @[fifo.scala 99:71]
  wire [135:0] fifo_banks_0_out = Look_up_table_read_first__io_out; // @[fifo.scala 42:{29,29}]
  wire [135:0] fifo_banks_1_out = Look_up_table_read_first__1_io_out; // @[fifo.scala 42:{29,29}]
  wire [135:0] _GEN_1 = 2'h1 == read_banks_points ? fifo_banks_1_out : fifo_banks_0_out; // @[fifo.scala 103:{30,30}]
  wire [135:0] fifo_banks_2_out = Look_up_table_read_first__2_io_out; // @[fifo.scala 42:{29,29}]
  wire [135:0] _GEN_2 = 2'h2 == read_banks_points ? fifo_banks_2_out : _GEN_1; // @[fifo.scala 103:{30,30}]
  wire [135:0] fifo_banks_3_out = Look_up_table_read_first__3_io_out; // @[fifo.scala 42:{29,29}]
  wire [135:0] _GEN_3 = 2'h3 == read_banks_points ? fifo_banks_3_out : _GEN_2; // @[fifo.scala 103:{30,30}]
  wire  _io_empty_T_1 = write_length_points == read_length_points; // @[fifo.scala 110:81]
  wire [2:0] _io_full_T_3 = _write_length_points_T_5 + 3'h1; // @[fifo.scala 112:98]
  wire [3:0] _io_full_T_7 = write_length_points + 4'h1; // @[fifo.scala 113:33]
  wire  _io_full_T_12 = _io_full_T_7 == read_length_points & (_fifo_banks_3_write_T_1 & read_banks_points == 2'h0); // @[fifo.scala 113:12]
  Look_up_table_read_first_ Look_up_table_read_first_ ( // @[fifo.scala 42:55]
    .clock(Look_up_table_read_first__clock),
    .reset(Look_up_table_read_first__reset),
    .io_ar_addr(Look_up_table_read_first__io_ar_addr),
    .io_aw_addr(Look_up_table_read_first__io_aw_addr),
    .io_write(Look_up_table_read_first__io_write),
    .io_in(Look_up_table_read_first__io_in),
    .io_out(Look_up_table_read_first__io_out)
  );
  Look_up_table_read_first_ Look_up_table_read_first__1 ( // @[fifo.scala 42:55]
    .clock(Look_up_table_read_first__1_clock),
    .reset(Look_up_table_read_first__1_reset),
    .io_ar_addr(Look_up_table_read_first__1_io_ar_addr),
    .io_aw_addr(Look_up_table_read_first__1_io_aw_addr),
    .io_write(Look_up_table_read_first__1_io_write),
    .io_in(Look_up_table_read_first__1_io_in),
    .io_out(Look_up_table_read_first__1_io_out)
  );
  Look_up_table_read_first_ Look_up_table_read_first__2 ( // @[fifo.scala 42:55]
    .clock(Look_up_table_read_first__2_clock),
    .reset(Look_up_table_read_first__2_reset),
    .io_ar_addr(Look_up_table_read_first__2_io_ar_addr),
    .io_aw_addr(Look_up_table_read_first__2_io_aw_addr),
    .io_write(Look_up_table_read_first__2_io_write),
    .io_in(Look_up_table_read_first__2_io_in),
    .io_out(Look_up_table_read_first__2_io_out)
  );
  Look_up_table_read_first_ Look_up_table_read_first__3 ( // @[fifo.scala 42:55]
    .clock(Look_up_table_read_first__3_clock),
    .reset(Look_up_table_read_first__3_reset),
    .io_ar_addr(Look_up_table_read_first__3_io_ar_addr),
    .io_aw_addr(Look_up_table_read_first__3_io_aw_addr),
    .io_write(Look_up_table_read_first__3_io_write),
    .io_in(Look_up_table_read_first__3_io_in),
    .io_out(Look_up_table_read_first__3_io_out)
  );
  assign io_read_out_0 = io_empty ? 136'h0 : _GEN_3; // @[fifo.scala 103:30]
  assign io_full = _io_empty_T_1 ? _io_full_T_3 == _read_length_points_T : _io_full_T_12; // @[fifo.scala 112:20]
  assign io_empty = write_banks_points == read_banks_points & write_length_points == read_length_points; // @[fifo.scala 110:58]
  assign Look_up_table_read_first__clock = clock;
  assign Look_up_table_read_first__reset = reset;
  assign Look_up_table_read_first__io_ar_addr = read_length_points; // @[fifo.scala 42:29 55:38]
  assign Look_up_table_read_first__io_aw_addr = write_length_points; // @[fifo.scala 42:29 50:38]
  assign Look_up_table_read_first__io_write = write_banks_points == 2'h0 & io_write_en[0]; // @[Mux.scala 81:58]
  assign Look_up_table_read_first__io_in = io_write_in_0; // @[fifo.scala 42:29 60:33]
  assign Look_up_table_read_first__1_clock = clock;
  assign Look_up_table_read_first__1_reset = reset;
  assign Look_up_table_read_first__1_io_ar_addr = read_length_points; // @[fifo.scala 42:29 55:38]
  assign Look_up_table_read_first__1_io_aw_addr = write_length_points; // @[fifo.scala 42:29 50:38]
  assign Look_up_table_read_first__1_io_write = write_banks_points == 2'h1 & io_write_en[0]; // @[Mux.scala 81:58]
  assign Look_up_table_read_first__1_io_in = io_write_in_0; // @[fifo.scala 42:29 60:33]
  assign Look_up_table_read_first__2_clock = clock;
  assign Look_up_table_read_first__2_reset = reset;
  assign Look_up_table_read_first__2_io_ar_addr = read_length_points; // @[fifo.scala 42:29 55:38]
  assign Look_up_table_read_first__2_io_aw_addr = write_length_points; // @[fifo.scala 42:29 50:38]
  assign Look_up_table_read_first__2_io_write = write_banks_points == 2'h2 & io_write_en[0]; // @[Mux.scala 81:58]
  assign Look_up_table_read_first__2_io_in = io_write_in_0; // @[fifo.scala 42:29 60:33]
  assign Look_up_table_read_first__3_clock = clock;
  assign Look_up_table_read_first__3_reset = reset;
  assign Look_up_table_read_first__3_io_ar_addr = read_length_points; // @[fifo.scala 42:29 55:38]
  assign Look_up_table_read_first__3_io_aw_addr = write_length_points; // @[fifo.scala 42:29 50:38]
  assign Look_up_table_read_first__3_io_write = write_banks_points == 2'h3 & io_write_en[0]; // @[Mux.scala 81:58]
  assign Look_up_table_read_first__3_io_in = io_write_in_0; // @[fifo.scala 42:29 60:33]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[fifo.scala 93:30]
      write_banks_points <= 2'h0;
    end else if (io_point_flush) begin // @[fifo.scala 93:53]
      write_banks_points <= 2'h0;
    end else if (point_write_tag) begin
      write_banks_points <= _write_banks_points_T_2;
    end else begin
      write_banks_points <= _write_banks_points_T_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[fifo.scala 97:31]
      write_length_points <= 4'h0;
    end else if (io_point_flush) begin // @[fifo.scala 97:54]
      write_length_points <= 4'h0;
    end else if (point_write_tag) begin
      write_length_points <= _write_length_points_T_4;
    end else begin
      write_length_points <= _write_length_points_T_11;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[fifo.scala 98:29]
      read_banks_points <= 2'h0;
    end else if (io_point_flush) begin
      read_banks_points <= 2'h0;
    end else begin
      read_banks_points <= _read_banks_points_T_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[fifo.scala 99:30]
      read_length_points <= 4'h0;
    end else if (io_point_flush) begin
      read_length_points <= 4'h0;
    end else begin
      read_length_points <= _read_length_points_T_6;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  write_banks_points = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  write_length_points = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  read_banks_points = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  read_length_points = _RAND_3[3:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    write_banks_points = 2'h0;
  end
  if (reset) begin
    write_length_points = 4'h0;
  end
  if (reset) begin
    read_banks_points = 2'h0;
  end
  if (reset) begin
    read_length_points = 4'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module pc_detail(
  input         clock,
  input         reset,
  input         io_stall,
  input         io_flush,
  input  [31:0] io_in_pc_value_in,
  output [31:0] io_out_pc_value_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] pc_value; // @[myCPU.scala 307:25]
  assign io_out_pc_value_out = pc_value; // @[myCPU.scala 310:25]
  always @(posedge clock) begin
    if (reset) begin // @[myCPU.scala 309:20]
      pc_value <= 32'hbfbffffc;
    end else if (io_flush) begin // @[myCPU.scala 309:60]
      pc_value <= 32'h0;
    end else if (io_stall) begin // @[myCPU.scala 309:77]
      pc_value <= io_in_pc_value_in;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc_value = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module pht_data_with_block_ram(
  input        clock,
  input        io_wen,
  input  [4:0] io_raddr,
  input  [4:0] io_waddr,
  input  [7:0] io_wdata,
  output [7:0] io_rdata
);
  wire  btb_data_ram_0_clka; // @[PHTS.scala 176:32]
  wire  btb_data_ram_0_clkb; // @[PHTS.scala 176:32]
  wire  btb_data_ram_0_ena; // @[PHTS.scala 176:32]
  wire  btb_data_ram_0_enb; // @[PHTS.scala 176:32]
  wire  btb_data_ram_0_wea; // @[PHTS.scala 176:32]
  wire [4:0] btb_data_ram_0_addra; // @[PHTS.scala 176:32]
  wire [7:0] btb_data_ram_0_dina; // @[PHTS.scala 176:32]
  wire [4:0] btb_data_ram_0_addrb; // @[PHTS.scala 176:32]
  wire [7:0] btb_data_ram_0_doutb; // @[PHTS.scala 176:32]
  pht_data_ram btb_data_ram_0 ( // @[PHTS.scala 176:32]
    .clka(btb_data_ram_0_clka),
    .clkb(btb_data_ram_0_clkb),
    .ena(btb_data_ram_0_ena),
    .enb(btb_data_ram_0_enb),
    .wea(btb_data_ram_0_wea),
    .addra(btb_data_ram_0_addra),
    .dina(btb_data_ram_0_dina),
    .addrb(btb_data_ram_0_addrb),
    .doutb(btb_data_ram_0_doutb)
  );
  assign io_rdata = btb_data_ram_0_doutb; // @[PHTS.scala 185:18]
  assign btb_data_ram_0_clka = clock; // @[PHTS.scala 177:37]
  assign btb_data_ram_0_clkb = clock; // @[PHTS.scala 178:37]
  assign btb_data_ram_0_ena = 1'h1; // @[PHTS.scala 179:29]
  assign btb_data_ram_0_enb = 1'h1; // @[PHTS.scala 180:29]
  assign btb_data_ram_0_wea = io_wen; // @[PHTS.scala 181:28]
  assign btb_data_ram_0_addra = io_waddr; // @[PHTS.scala 182:29]
  assign btb_data_ram_0_dina = io_wdata; // @[PHTS.scala 184:28]
  assign btb_data_ram_0_addrb = io_raddr; // @[PHTS.scala 183:29]
endmodule
module PHTS_with_block_ram(
  input        clock,
  input        reset,
  input  [6:0] io_ar_addr,
  input  [2:0] io_ar_pht_addr,
  input  [6:0] io_aw_addr,
  input  [2:0] io_aw_pht_addr,
  input        io_write,
  input  [7:0] io_in,
  output [7:0] io_pht_out,
  output [1:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  pht_data_with_block_ram_clock; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_io_wen; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_io_raddr; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_io_waddr; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_io_wdata; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_io_rdata; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_1_clock; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_1_io_wen; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_1_io_raddr; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_1_io_waddr; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_1_io_wdata; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_1_io_rdata; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_2_clock; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_2_io_wen; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_2_io_raddr; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_2_io_waddr; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_2_io_wdata; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_2_io_rdata; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_3_clock; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_3_io_wen; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_3_io_raddr; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_3_io_waddr; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_3_io_wdata; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_3_io_rdata; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_4_clock; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_4_io_wen; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_4_io_raddr; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_4_io_waddr; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_4_io_wdata; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_4_io_rdata; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_5_clock; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_5_io_wen; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_5_io_raddr; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_5_io_waddr; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_5_io_wdata; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_5_io_rdata; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_6_clock; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_6_io_wen; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_6_io_raddr; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_6_io_waddr; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_6_io_wdata; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_6_io_rdata; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_7_clock; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_7_io_wen; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_7_io_raddr; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_7_io_waddr; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_7_io_wdata; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_7_io_rdata; // @[PHTS.scala 205:45]
  reg [6:0] raddr_reg; // @[PHTS.scala 213:28]
  reg [7:0] ways_araddr_reg; // @[PHTS.scala 214:34]
  wire [7:0] phts_0_rdata = pht_data_with_block_ram_io_rdata; // @[PHTS.scala 205:{23,23}]
  wire [7:0] phts_1_rdata = pht_data_with_block_ram_1_io_rdata; // @[PHTS.scala 205:{23,23}]
  wire [7:0] _GEN_1 = 3'h1 == ways_araddr_reg[2:0] ? phts_1_rdata : phts_0_rdata; // @[PHTS.scala 217:{67,67}]
  wire [7:0] phts_2_rdata = pht_data_with_block_ram_2_io_rdata; // @[PHTS.scala 205:{23,23}]
  wire [7:0] _GEN_2 = 3'h2 == ways_araddr_reg[2:0] ? phts_2_rdata : _GEN_1; // @[PHTS.scala 217:{67,67}]
  wire [7:0] phts_3_rdata = pht_data_with_block_ram_3_io_rdata; // @[PHTS.scala 205:{23,23}]
  wire [7:0] _GEN_3 = 3'h3 == ways_araddr_reg[2:0] ? phts_3_rdata : _GEN_2; // @[PHTS.scala 217:{67,67}]
  wire [7:0] phts_4_rdata = pht_data_with_block_ram_4_io_rdata; // @[PHTS.scala 205:{23,23}]
  wire [7:0] _GEN_4 = 3'h4 == ways_araddr_reg[2:0] ? phts_4_rdata : _GEN_3; // @[PHTS.scala 217:{67,67}]
  wire [7:0] phts_5_rdata = pht_data_with_block_ram_5_io_rdata; // @[PHTS.scala 205:{23,23}]
  wire [7:0] _GEN_5 = 3'h5 == ways_araddr_reg[2:0] ? phts_5_rdata : _GEN_4; // @[PHTS.scala 217:{67,67}]
  wire [7:0] phts_6_rdata = pht_data_with_block_ram_6_io_rdata; // @[PHTS.scala 205:{23,23}]
  wire [7:0] _GEN_6 = 3'h6 == ways_araddr_reg[2:0] ? phts_6_rdata : _GEN_5; // @[PHTS.scala 217:{67,67}]
  wire [7:0] phts_7_rdata = pht_data_with_block_ram_7_io_rdata; // @[PHTS.scala 205:{23,23}]
  wire [7:0] _GEN_7 = 3'h7 == ways_araddr_reg[2:0] ? phts_7_rdata : _GEN_6; // @[PHTS.scala 217:{67,67}]
  wire [1:0] _io_out_T_10 = 2'h0 == raddr_reg[1:0] ? _GEN_7[1:0] : _GEN_7[7:6]; // @[Mux.scala 81:58]
  wire [1:0] _io_out_T_12 = 2'h1 == raddr_reg[1:0] ? _GEN_7[3:2] : _io_out_T_10; // @[Mux.scala 81:58]
  pht_data_with_block_ram pht_data_with_block_ram ( // @[PHTS.scala 205:45]
    .clock(pht_data_with_block_ram_clock),
    .io_wen(pht_data_with_block_ram_io_wen),
    .io_raddr(pht_data_with_block_ram_io_raddr),
    .io_waddr(pht_data_with_block_ram_io_waddr),
    .io_wdata(pht_data_with_block_ram_io_wdata),
    .io_rdata(pht_data_with_block_ram_io_rdata)
  );
  pht_data_with_block_ram pht_data_with_block_ram_1 ( // @[PHTS.scala 205:45]
    .clock(pht_data_with_block_ram_1_clock),
    .io_wen(pht_data_with_block_ram_1_io_wen),
    .io_raddr(pht_data_with_block_ram_1_io_raddr),
    .io_waddr(pht_data_with_block_ram_1_io_waddr),
    .io_wdata(pht_data_with_block_ram_1_io_wdata),
    .io_rdata(pht_data_with_block_ram_1_io_rdata)
  );
  pht_data_with_block_ram pht_data_with_block_ram_2 ( // @[PHTS.scala 205:45]
    .clock(pht_data_with_block_ram_2_clock),
    .io_wen(pht_data_with_block_ram_2_io_wen),
    .io_raddr(pht_data_with_block_ram_2_io_raddr),
    .io_waddr(pht_data_with_block_ram_2_io_waddr),
    .io_wdata(pht_data_with_block_ram_2_io_wdata),
    .io_rdata(pht_data_with_block_ram_2_io_rdata)
  );
  pht_data_with_block_ram pht_data_with_block_ram_3 ( // @[PHTS.scala 205:45]
    .clock(pht_data_with_block_ram_3_clock),
    .io_wen(pht_data_with_block_ram_3_io_wen),
    .io_raddr(pht_data_with_block_ram_3_io_raddr),
    .io_waddr(pht_data_with_block_ram_3_io_waddr),
    .io_wdata(pht_data_with_block_ram_3_io_wdata),
    .io_rdata(pht_data_with_block_ram_3_io_rdata)
  );
  pht_data_with_block_ram pht_data_with_block_ram_4 ( // @[PHTS.scala 205:45]
    .clock(pht_data_with_block_ram_4_clock),
    .io_wen(pht_data_with_block_ram_4_io_wen),
    .io_raddr(pht_data_with_block_ram_4_io_raddr),
    .io_waddr(pht_data_with_block_ram_4_io_waddr),
    .io_wdata(pht_data_with_block_ram_4_io_wdata),
    .io_rdata(pht_data_with_block_ram_4_io_rdata)
  );
  pht_data_with_block_ram pht_data_with_block_ram_5 ( // @[PHTS.scala 205:45]
    .clock(pht_data_with_block_ram_5_clock),
    .io_wen(pht_data_with_block_ram_5_io_wen),
    .io_raddr(pht_data_with_block_ram_5_io_raddr),
    .io_waddr(pht_data_with_block_ram_5_io_waddr),
    .io_wdata(pht_data_with_block_ram_5_io_wdata),
    .io_rdata(pht_data_with_block_ram_5_io_rdata)
  );
  pht_data_with_block_ram pht_data_with_block_ram_6 ( // @[PHTS.scala 205:45]
    .clock(pht_data_with_block_ram_6_clock),
    .io_wen(pht_data_with_block_ram_6_io_wen),
    .io_raddr(pht_data_with_block_ram_6_io_raddr),
    .io_waddr(pht_data_with_block_ram_6_io_waddr),
    .io_wdata(pht_data_with_block_ram_6_io_wdata),
    .io_rdata(pht_data_with_block_ram_6_io_rdata)
  );
  pht_data_with_block_ram pht_data_with_block_ram_7 ( // @[PHTS.scala 205:45]
    .clock(pht_data_with_block_ram_7_clock),
    .io_wen(pht_data_with_block_ram_7_io_wen),
    .io_raddr(pht_data_with_block_ram_7_io_raddr),
    .io_waddr(pht_data_with_block_ram_7_io_waddr),
    .io_wdata(pht_data_with_block_ram_7_io_wdata),
    .io_rdata(pht_data_with_block_ram_7_io_rdata)
  );
  assign io_pht_out = 3'h7 == ways_araddr_reg[2:0] ? phts_7_rdata : _GEN_6; // @[PHTS.scala 222:{16,16}]
  assign io_out = 2'h2 == raddr_reg[1:0] ? _GEN_7[5:4] : _io_out_T_12; // @[Mux.scala 81:58]
  assign pht_data_with_block_ram_clock = clock;
  assign pht_data_with_block_ram_io_wen = io_aw_pht_addr == 3'h0 & io_write; // @[PHTS.scala 207:52]
  assign pht_data_with_block_ram_io_raddr = io_ar_addr[6:2]; // @[PHTS.scala 210:36]
  assign pht_data_with_block_ram_io_waddr = io_aw_addr[6:2]; // @[PHTS.scala 211:36]
  assign pht_data_with_block_ram_io_wdata = io_in; // @[PHTS.scala 205:23 209:23]
  assign pht_data_with_block_ram_1_clock = clock;
  assign pht_data_with_block_ram_1_io_wen = io_aw_pht_addr == 3'h1 & io_write; // @[PHTS.scala 207:52]
  assign pht_data_with_block_ram_1_io_raddr = io_ar_addr[6:2]; // @[PHTS.scala 210:36]
  assign pht_data_with_block_ram_1_io_waddr = io_aw_addr[6:2]; // @[PHTS.scala 211:36]
  assign pht_data_with_block_ram_1_io_wdata = io_in; // @[PHTS.scala 205:23 209:23]
  assign pht_data_with_block_ram_2_clock = clock;
  assign pht_data_with_block_ram_2_io_wen = io_aw_pht_addr == 3'h2 & io_write; // @[PHTS.scala 207:52]
  assign pht_data_with_block_ram_2_io_raddr = io_ar_addr[6:2]; // @[PHTS.scala 210:36]
  assign pht_data_with_block_ram_2_io_waddr = io_aw_addr[6:2]; // @[PHTS.scala 211:36]
  assign pht_data_with_block_ram_2_io_wdata = io_in; // @[PHTS.scala 205:23 209:23]
  assign pht_data_with_block_ram_3_clock = clock;
  assign pht_data_with_block_ram_3_io_wen = io_aw_pht_addr == 3'h3 & io_write; // @[PHTS.scala 207:52]
  assign pht_data_with_block_ram_3_io_raddr = io_ar_addr[6:2]; // @[PHTS.scala 210:36]
  assign pht_data_with_block_ram_3_io_waddr = io_aw_addr[6:2]; // @[PHTS.scala 211:36]
  assign pht_data_with_block_ram_3_io_wdata = io_in; // @[PHTS.scala 205:23 209:23]
  assign pht_data_with_block_ram_4_clock = clock;
  assign pht_data_with_block_ram_4_io_wen = io_aw_pht_addr == 3'h4 & io_write; // @[PHTS.scala 207:52]
  assign pht_data_with_block_ram_4_io_raddr = io_ar_addr[6:2]; // @[PHTS.scala 210:36]
  assign pht_data_with_block_ram_4_io_waddr = io_aw_addr[6:2]; // @[PHTS.scala 211:36]
  assign pht_data_with_block_ram_4_io_wdata = io_in; // @[PHTS.scala 205:23 209:23]
  assign pht_data_with_block_ram_5_clock = clock;
  assign pht_data_with_block_ram_5_io_wen = io_aw_pht_addr == 3'h5 & io_write; // @[PHTS.scala 207:52]
  assign pht_data_with_block_ram_5_io_raddr = io_ar_addr[6:2]; // @[PHTS.scala 210:36]
  assign pht_data_with_block_ram_5_io_waddr = io_aw_addr[6:2]; // @[PHTS.scala 211:36]
  assign pht_data_with_block_ram_5_io_wdata = io_in; // @[PHTS.scala 205:23 209:23]
  assign pht_data_with_block_ram_6_clock = clock;
  assign pht_data_with_block_ram_6_io_wen = io_aw_pht_addr == 3'h6 & io_write; // @[PHTS.scala 207:52]
  assign pht_data_with_block_ram_6_io_raddr = io_ar_addr[6:2]; // @[PHTS.scala 210:36]
  assign pht_data_with_block_ram_6_io_waddr = io_aw_addr[6:2]; // @[PHTS.scala 211:36]
  assign pht_data_with_block_ram_6_io_wdata = io_in; // @[PHTS.scala 205:23 209:23]
  assign pht_data_with_block_ram_7_clock = clock;
  assign pht_data_with_block_ram_7_io_wen = io_aw_pht_addr == 3'h7 & io_write; // @[PHTS.scala 207:52]
  assign pht_data_with_block_ram_7_io_raddr = io_ar_addr[6:2]; // @[PHTS.scala 210:36]
  assign pht_data_with_block_ram_7_io_waddr = io_aw_addr[6:2]; // @[PHTS.scala 211:36]
  assign pht_data_with_block_ram_7_io_wdata = io_in; // @[PHTS.scala 205:23 209:23]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PHTS.scala 213:28]
      raddr_reg <= 7'h0; // @[PHTS.scala 213:28]
    end else begin
      raddr_reg <= io_ar_addr; // @[PHTS.scala 215:15]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PHTS.scala 214:34]
      ways_araddr_reg <= 8'h0; // @[PHTS.scala 214:34]
    end else begin
      ways_araddr_reg <= {{5'd0}, io_ar_pht_addr}; // @[PHTS.scala 216:21]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  raddr_reg = _RAND_0[6:0];
  _RAND_1 = {1{`RANDOM}};
  ways_araddr_reg = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    raddr_reg = 7'h0;
  end
  if (reset) begin
    ways_araddr_reg = 8'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PHTS_banks_oneissue_block_ram(
  input        clock,
  input        reset,
  input  [1:0] io_ar_bank_sel,
  input  [6:0] io_ar_addr_L,
  input  [2:0] io_ar_pht_addr,
  input  [6:0] io_aw_addr,
  input  [2:0] io_aw_pht_addr,
  input  [1:0] io_aw_bank_sel,
  input        io_write,
  input  [7:0] io_in,
  output [1:0] io_out_L,
  output [7:0] io_pht_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  PHTS_with_block_ram_clock; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_reset; // @[PHTS.scala 250:55]
  wire [6:0] PHTS_with_block_ram_io_ar_addr; // @[PHTS.scala 250:55]
  wire [2:0] PHTS_with_block_ram_io_ar_pht_addr; // @[PHTS.scala 250:55]
  wire [6:0] PHTS_with_block_ram_io_aw_addr; // @[PHTS.scala 250:55]
  wire [2:0] PHTS_with_block_ram_io_aw_pht_addr; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_io_write; // @[PHTS.scala 250:55]
  wire [7:0] PHTS_with_block_ram_io_in; // @[PHTS.scala 250:55]
  wire [7:0] PHTS_with_block_ram_io_pht_out; // @[PHTS.scala 250:55]
  wire [1:0] PHTS_with_block_ram_io_out; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_1_clock; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_1_reset; // @[PHTS.scala 250:55]
  wire [6:0] PHTS_with_block_ram_1_io_ar_addr; // @[PHTS.scala 250:55]
  wire [2:0] PHTS_with_block_ram_1_io_ar_pht_addr; // @[PHTS.scala 250:55]
  wire [6:0] PHTS_with_block_ram_1_io_aw_addr; // @[PHTS.scala 250:55]
  wire [2:0] PHTS_with_block_ram_1_io_aw_pht_addr; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_1_io_write; // @[PHTS.scala 250:55]
  wire [7:0] PHTS_with_block_ram_1_io_in; // @[PHTS.scala 250:55]
  wire [7:0] PHTS_with_block_ram_1_io_pht_out; // @[PHTS.scala 250:55]
  wire [1:0] PHTS_with_block_ram_1_io_out; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_2_clock; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_2_reset; // @[PHTS.scala 250:55]
  wire [6:0] PHTS_with_block_ram_2_io_ar_addr; // @[PHTS.scala 250:55]
  wire [2:0] PHTS_with_block_ram_2_io_ar_pht_addr; // @[PHTS.scala 250:55]
  wire [6:0] PHTS_with_block_ram_2_io_aw_addr; // @[PHTS.scala 250:55]
  wire [2:0] PHTS_with_block_ram_2_io_aw_pht_addr; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_2_io_write; // @[PHTS.scala 250:55]
  wire [7:0] PHTS_with_block_ram_2_io_in; // @[PHTS.scala 250:55]
  wire [7:0] PHTS_with_block_ram_2_io_pht_out; // @[PHTS.scala 250:55]
  wire [1:0] PHTS_with_block_ram_2_io_out; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_3_clock; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_3_reset; // @[PHTS.scala 250:55]
  wire [6:0] PHTS_with_block_ram_3_io_ar_addr; // @[PHTS.scala 250:55]
  wire [2:0] PHTS_with_block_ram_3_io_ar_pht_addr; // @[PHTS.scala 250:55]
  wire [6:0] PHTS_with_block_ram_3_io_aw_addr; // @[PHTS.scala 250:55]
  wire [2:0] PHTS_with_block_ram_3_io_aw_pht_addr; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_3_io_write; // @[PHTS.scala 250:55]
  wire [7:0] PHTS_with_block_ram_3_io_in; // @[PHTS.scala 250:55]
  wire [7:0] PHTS_with_block_ram_3_io_pht_out; // @[PHTS.scala 250:55]
  wire [1:0] PHTS_with_block_ram_3_io_out; // @[PHTS.scala 250:55]
  reg [1:0] ar_bank_sel_reg; // @[PHTS.scala 261:34]
  wire [1:0] phts_banks_0_out = PHTS_with_block_ram_io_out; // @[PHTS.scala 250:{29,29}]
  wire [1:0] phts_banks_1_out = PHTS_with_block_ram_1_io_out; // @[PHTS.scala 250:{29,29}]
  wire [1:0] _GEN_1 = 2'h1 == ar_bank_sel_reg ? phts_banks_1_out : phts_banks_0_out; // @[PHTS.scala 263:{14,14}]
  wire [1:0] phts_banks_2_out = PHTS_with_block_ram_2_io_out; // @[PHTS.scala 250:{29,29}]
  wire [1:0] _GEN_2 = 2'h2 == ar_bank_sel_reg ? phts_banks_2_out : _GEN_1; // @[PHTS.scala 263:{14,14}]
  wire [1:0] phts_banks_3_out = PHTS_with_block_ram_3_io_out; // @[PHTS.scala 250:{29,29}]
  wire [7:0] phts_banks_0_pht_out = PHTS_with_block_ram_io_pht_out; // @[PHTS.scala 250:{29,29}]
  wire [7:0] phts_banks_1_pht_out = PHTS_with_block_ram_1_io_pht_out; // @[PHTS.scala 250:{29,29}]
  wire [7:0] _GEN_5 = 2'h1 == ar_bank_sel_reg ? phts_banks_1_pht_out : phts_banks_0_pht_out; // @[PHTS.scala 266:{16,16}]
  wire [7:0] phts_banks_2_pht_out = PHTS_with_block_ram_2_io_pht_out; // @[PHTS.scala 250:{29,29}]
  wire [7:0] _GEN_6 = 2'h2 == ar_bank_sel_reg ? phts_banks_2_pht_out : _GEN_5; // @[PHTS.scala 266:{16,16}]
  wire [7:0] phts_banks_3_pht_out = PHTS_with_block_ram_3_io_pht_out; // @[PHTS.scala 250:{29,29}]
  PHTS_with_block_ram PHTS_with_block_ram ( // @[PHTS.scala 250:55]
    .clock(PHTS_with_block_ram_clock),
    .reset(PHTS_with_block_ram_reset),
    .io_ar_addr(PHTS_with_block_ram_io_ar_addr),
    .io_ar_pht_addr(PHTS_with_block_ram_io_ar_pht_addr),
    .io_aw_addr(PHTS_with_block_ram_io_aw_addr),
    .io_aw_pht_addr(PHTS_with_block_ram_io_aw_pht_addr),
    .io_write(PHTS_with_block_ram_io_write),
    .io_in(PHTS_with_block_ram_io_in),
    .io_pht_out(PHTS_with_block_ram_io_pht_out),
    .io_out(PHTS_with_block_ram_io_out)
  );
  PHTS_with_block_ram PHTS_with_block_ram_1 ( // @[PHTS.scala 250:55]
    .clock(PHTS_with_block_ram_1_clock),
    .reset(PHTS_with_block_ram_1_reset),
    .io_ar_addr(PHTS_with_block_ram_1_io_ar_addr),
    .io_ar_pht_addr(PHTS_with_block_ram_1_io_ar_pht_addr),
    .io_aw_addr(PHTS_with_block_ram_1_io_aw_addr),
    .io_aw_pht_addr(PHTS_with_block_ram_1_io_aw_pht_addr),
    .io_write(PHTS_with_block_ram_1_io_write),
    .io_in(PHTS_with_block_ram_1_io_in),
    .io_pht_out(PHTS_with_block_ram_1_io_pht_out),
    .io_out(PHTS_with_block_ram_1_io_out)
  );
  PHTS_with_block_ram PHTS_with_block_ram_2 ( // @[PHTS.scala 250:55]
    .clock(PHTS_with_block_ram_2_clock),
    .reset(PHTS_with_block_ram_2_reset),
    .io_ar_addr(PHTS_with_block_ram_2_io_ar_addr),
    .io_ar_pht_addr(PHTS_with_block_ram_2_io_ar_pht_addr),
    .io_aw_addr(PHTS_with_block_ram_2_io_aw_addr),
    .io_aw_pht_addr(PHTS_with_block_ram_2_io_aw_pht_addr),
    .io_write(PHTS_with_block_ram_2_io_write),
    .io_in(PHTS_with_block_ram_2_io_in),
    .io_pht_out(PHTS_with_block_ram_2_io_pht_out),
    .io_out(PHTS_with_block_ram_2_io_out)
  );
  PHTS_with_block_ram PHTS_with_block_ram_3 ( // @[PHTS.scala 250:55]
    .clock(PHTS_with_block_ram_3_clock),
    .reset(PHTS_with_block_ram_3_reset),
    .io_ar_addr(PHTS_with_block_ram_3_io_ar_addr),
    .io_ar_pht_addr(PHTS_with_block_ram_3_io_ar_pht_addr),
    .io_aw_addr(PHTS_with_block_ram_3_io_aw_addr),
    .io_aw_pht_addr(PHTS_with_block_ram_3_io_aw_pht_addr),
    .io_write(PHTS_with_block_ram_3_io_write),
    .io_in(PHTS_with_block_ram_3_io_in),
    .io_pht_out(PHTS_with_block_ram_3_io_pht_out),
    .io_out(PHTS_with_block_ram_3_io_out)
  );
  assign io_out_L = 2'h3 == ar_bank_sel_reg ? phts_banks_3_out : _GEN_2; // @[PHTS.scala 263:{14,14}]
  assign io_pht_out = 2'h3 == ar_bank_sel_reg ? phts_banks_3_pht_out : _GEN_6; // @[PHTS.scala 266:{16,16}]
  assign PHTS_with_block_ram_clock = clock;
  assign PHTS_with_block_ram_reset = reset;
  assign PHTS_with_block_ram_io_ar_addr = io_ar_addr_L; // @[PHTS.scala 250:29 254:31]
  assign PHTS_with_block_ram_io_ar_pht_addr = io_ar_pht_addr; // @[PHTS.scala 250:29 257:35]
  assign PHTS_with_block_ram_io_aw_addr = io_aw_addr; // @[PHTS.scala 250:29 258:31]
  assign PHTS_with_block_ram_io_aw_pht_addr = io_aw_pht_addr; // @[PHTS.scala 250:29 259:35]
  assign PHTS_with_block_ram_io_write = io_aw_bank_sel == 2'h0 & io_write; // @[PHTS.scala 252:60]
  assign PHTS_with_block_ram_io_in = io_in; // @[PHTS.scala 250:29 253:26]
  assign PHTS_with_block_ram_1_clock = clock;
  assign PHTS_with_block_ram_1_reset = reset;
  assign PHTS_with_block_ram_1_io_ar_addr = io_ar_addr_L; // @[PHTS.scala 250:29 254:31]
  assign PHTS_with_block_ram_1_io_ar_pht_addr = io_ar_pht_addr; // @[PHTS.scala 250:29 257:35]
  assign PHTS_with_block_ram_1_io_aw_addr = io_aw_addr; // @[PHTS.scala 250:29 258:31]
  assign PHTS_with_block_ram_1_io_aw_pht_addr = io_aw_pht_addr; // @[PHTS.scala 250:29 259:35]
  assign PHTS_with_block_ram_1_io_write = io_aw_bank_sel == 2'h1 & io_write; // @[PHTS.scala 252:60]
  assign PHTS_with_block_ram_1_io_in = io_in; // @[PHTS.scala 250:29 253:26]
  assign PHTS_with_block_ram_2_clock = clock;
  assign PHTS_with_block_ram_2_reset = reset;
  assign PHTS_with_block_ram_2_io_ar_addr = io_ar_addr_L; // @[PHTS.scala 250:29 254:31]
  assign PHTS_with_block_ram_2_io_ar_pht_addr = io_ar_pht_addr; // @[PHTS.scala 250:29 257:35]
  assign PHTS_with_block_ram_2_io_aw_addr = io_aw_addr; // @[PHTS.scala 250:29 258:31]
  assign PHTS_with_block_ram_2_io_aw_pht_addr = io_aw_pht_addr; // @[PHTS.scala 250:29 259:35]
  assign PHTS_with_block_ram_2_io_write = io_aw_bank_sel == 2'h2 & io_write; // @[PHTS.scala 252:60]
  assign PHTS_with_block_ram_2_io_in = io_in; // @[PHTS.scala 250:29 253:26]
  assign PHTS_with_block_ram_3_clock = clock;
  assign PHTS_with_block_ram_3_reset = reset;
  assign PHTS_with_block_ram_3_io_ar_addr = io_ar_addr_L; // @[PHTS.scala 250:29 254:31]
  assign PHTS_with_block_ram_3_io_ar_pht_addr = io_ar_pht_addr; // @[PHTS.scala 250:29 257:35]
  assign PHTS_with_block_ram_3_io_aw_addr = io_aw_addr; // @[PHTS.scala 250:29 258:31]
  assign PHTS_with_block_ram_3_io_aw_pht_addr = io_aw_pht_addr; // @[PHTS.scala 250:29 259:35]
  assign PHTS_with_block_ram_3_io_write = io_aw_bank_sel == 2'h3 & io_write; // @[PHTS.scala 252:60]
  assign PHTS_with_block_ram_3_io_in = io_in; // @[PHTS.scala 250:29 253:26]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PHTS.scala 261:34]
      ar_bank_sel_reg <= 2'h0; // @[PHTS.scala 261:34]
    end else begin
      ar_bank_sel_reg <= io_ar_bank_sel; // @[PHTS.scala 262:21]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ar_bank_sel_reg = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    ar_bank_sel_reg = 2'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BHT(
  input        clock,
  input        reset,
  input  [6:0] io_ar_addr,
  input  [6:0] io_aw_addr,
  input        io_write,
  input  [2:0] io_in,
  output [2:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] bht_0; // @[BHT.scala 20:22]
  reg [2:0] bht_1; // @[BHT.scala 20:22]
  reg [2:0] bht_2; // @[BHT.scala 20:22]
  reg [2:0] bht_3; // @[BHT.scala 20:22]
  reg [2:0] bht_4; // @[BHT.scala 20:22]
  reg [2:0] bht_5; // @[BHT.scala 20:22]
  reg [2:0] bht_6; // @[BHT.scala 20:22]
  reg [2:0] bht_7; // @[BHT.scala 20:22]
  reg [2:0] bht_8; // @[BHT.scala 20:22]
  reg [2:0] bht_9; // @[BHT.scala 20:22]
  reg [2:0] bht_10; // @[BHT.scala 20:22]
  reg [2:0] bht_11; // @[BHT.scala 20:22]
  reg [2:0] bht_12; // @[BHT.scala 20:22]
  reg [2:0] bht_13; // @[BHT.scala 20:22]
  reg [2:0] bht_14; // @[BHT.scala 20:22]
  reg [2:0] bht_15; // @[BHT.scala 20:22]
  reg [2:0] bht_16; // @[BHT.scala 20:22]
  reg [2:0] bht_17; // @[BHT.scala 20:22]
  reg [2:0] bht_18; // @[BHT.scala 20:22]
  reg [2:0] bht_19; // @[BHT.scala 20:22]
  reg [2:0] bht_20; // @[BHT.scala 20:22]
  reg [2:0] bht_21; // @[BHT.scala 20:22]
  reg [2:0] bht_22; // @[BHT.scala 20:22]
  reg [2:0] bht_23; // @[BHT.scala 20:22]
  reg [2:0] bht_24; // @[BHT.scala 20:22]
  reg [2:0] bht_25; // @[BHT.scala 20:22]
  reg [2:0] bht_26; // @[BHT.scala 20:22]
  reg [2:0] bht_27; // @[BHT.scala 20:22]
  reg [2:0] bht_28; // @[BHT.scala 20:22]
  reg [2:0] bht_29; // @[BHT.scala 20:22]
  reg [2:0] bht_30; // @[BHT.scala 20:22]
  reg [2:0] bht_31; // @[BHT.scala 20:22]
  reg [2:0] bht_32; // @[BHT.scala 20:22]
  reg [2:0] bht_33; // @[BHT.scala 20:22]
  reg [2:0] bht_34; // @[BHT.scala 20:22]
  reg [2:0] bht_35; // @[BHT.scala 20:22]
  reg [2:0] bht_36; // @[BHT.scala 20:22]
  reg [2:0] bht_37; // @[BHT.scala 20:22]
  reg [2:0] bht_38; // @[BHT.scala 20:22]
  reg [2:0] bht_39; // @[BHT.scala 20:22]
  reg [2:0] bht_40; // @[BHT.scala 20:22]
  reg [2:0] bht_41; // @[BHT.scala 20:22]
  reg [2:0] bht_42; // @[BHT.scala 20:22]
  reg [2:0] bht_43; // @[BHT.scala 20:22]
  reg [2:0] bht_44; // @[BHT.scala 20:22]
  reg [2:0] bht_45; // @[BHT.scala 20:22]
  reg [2:0] bht_46; // @[BHT.scala 20:22]
  reg [2:0] bht_47; // @[BHT.scala 20:22]
  reg [2:0] bht_48; // @[BHT.scala 20:22]
  reg [2:0] bht_49; // @[BHT.scala 20:22]
  reg [2:0] bht_50; // @[BHT.scala 20:22]
  reg [2:0] bht_51; // @[BHT.scala 20:22]
  reg [2:0] bht_52; // @[BHT.scala 20:22]
  reg [2:0] bht_53; // @[BHT.scala 20:22]
  reg [2:0] bht_54; // @[BHT.scala 20:22]
  reg [2:0] bht_55; // @[BHT.scala 20:22]
  reg [2:0] bht_56; // @[BHT.scala 20:22]
  reg [2:0] bht_57; // @[BHT.scala 20:22]
  reg [2:0] bht_58; // @[BHT.scala 20:22]
  reg [2:0] bht_59; // @[BHT.scala 20:22]
  reg [2:0] bht_60; // @[BHT.scala 20:22]
  reg [2:0] bht_61; // @[BHT.scala 20:22]
  reg [2:0] bht_62; // @[BHT.scala 20:22]
  reg [2:0] bht_63; // @[BHT.scala 20:22]
  reg [2:0] bht_64; // @[BHT.scala 20:22]
  reg [2:0] bht_65; // @[BHT.scala 20:22]
  reg [2:0] bht_66; // @[BHT.scala 20:22]
  reg [2:0] bht_67; // @[BHT.scala 20:22]
  reg [2:0] bht_68; // @[BHT.scala 20:22]
  reg [2:0] bht_69; // @[BHT.scala 20:22]
  reg [2:0] bht_70; // @[BHT.scala 20:22]
  reg [2:0] bht_71; // @[BHT.scala 20:22]
  reg [2:0] bht_72; // @[BHT.scala 20:22]
  reg [2:0] bht_73; // @[BHT.scala 20:22]
  reg [2:0] bht_74; // @[BHT.scala 20:22]
  reg [2:0] bht_75; // @[BHT.scala 20:22]
  reg [2:0] bht_76; // @[BHT.scala 20:22]
  reg [2:0] bht_77; // @[BHT.scala 20:22]
  reg [2:0] bht_78; // @[BHT.scala 20:22]
  reg [2:0] bht_79; // @[BHT.scala 20:22]
  reg [2:0] bht_80; // @[BHT.scala 20:22]
  reg [2:0] bht_81; // @[BHT.scala 20:22]
  reg [2:0] bht_82; // @[BHT.scala 20:22]
  reg [2:0] bht_83; // @[BHT.scala 20:22]
  reg [2:0] bht_84; // @[BHT.scala 20:22]
  reg [2:0] bht_85; // @[BHT.scala 20:22]
  reg [2:0] bht_86; // @[BHT.scala 20:22]
  reg [2:0] bht_87; // @[BHT.scala 20:22]
  reg [2:0] bht_88; // @[BHT.scala 20:22]
  reg [2:0] bht_89; // @[BHT.scala 20:22]
  reg [2:0] bht_90; // @[BHT.scala 20:22]
  reg [2:0] bht_91; // @[BHT.scala 20:22]
  reg [2:0] bht_92; // @[BHT.scala 20:22]
  reg [2:0] bht_93; // @[BHT.scala 20:22]
  reg [2:0] bht_94; // @[BHT.scala 20:22]
  reg [2:0] bht_95; // @[BHT.scala 20:22]
  reg [2:0] bht_96; // @[BHT.scala 20:22]
  reg [2:0] bht_97; // @[BHT.scala 20:22]
  reg [2:0] bht_98; // @[BHT.scala 20:22]
  reg [2:0] bht_99; // @[BHT.scala 20:22]
  reg [2:0] bht_100; // @[BHT.scala 20:22]
  reg [2:0] bht_101; // @[BHT.scala 20:22]
  reg [2:0] bht_102; // @[BHT.scala 20:22]
  reg [2:0] bht_103; // @[BHT.scala 20:22]
  reg [2:0] bht_104; // @[BHT.scala 20:22]
  reg [2:0] bht_105; // @[BHT.scala 20:22]
  reg [2:0] bht_106; // @[BHT.scala 20:22]
  reg [2:0] bht_107; // @[BHT.scala 20:22]
  reg [2:0] bht_108; // @[BHT.scala 20:22]
  reg [2:0] bht_109; // @[BHT.scala 20:22]
  reg [2:0] bht_110; // @[BHT.scala 20:22]
  reg [2:0] bht_111; // @[BHT.scala 20:22]
  reg [2:0] bht_112; // @[BHT.scala 20:22]
  reg [2:0] bht_113; // @[BHT.scala 20:22]
  reg [2:0] bht_114; // @[BHT.scala 20:22]
  reg [2:0] bht_115; // @[BHT.scala 20:22]
  reg [2:0] bht_116; // @[BHT.scala 20:22]
  reg [2:0] bht_117; // @[BHT.scala 20:22]
  reg [2:0] bht_118; // @[BHT.scala 20:22]
  reg [2:0] bht_119; // @[BHT.scala 20:22]
  reg [2:0] bht_120; // @[BHT.scala 20:22]
  reg [2:0] bht_121; // @[BHT.scala 20:22]
  reg [2:0] bht_122; // @[BHT.scala 20:22]
  reg [2:0] bht_123; // @[BHT.scala 20:22]
  reg [2:0] bht_124; // @[BHT.scala 20:22]
  reg [2:0] bht_125; // @[BHT.scala 20:22]
  reg [2:0] bht_126; // @[BHT.scala 20:22]
  reg [2:0] bht_127; // @[BHT.scala 20:22]
  wire [2:0] _GEN_1 = 7'h1 == io_ar_addr ? bht_1 : bht_0; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_2 = 7'h2 == io_ar_addr ? bht_2 : _GEN_1; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_3 = 7'h3 == io_ar_addr ? bht_3 : _GEN_2; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_4 = 7'h4 == io_ar_addr ? bht_4 : _GEN_3; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_5 = 7'h5 == io_ar_addr ? bht_5 : _GEN_4; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_6 = 7'h6 == io_ar_addr ? bht_6 : _GEN_5; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_7 = 7'h7 == io_ar_addr ? bht_7 : _GEN_6; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_8 = 7'h8 == io_ar_addr ? bht_8 : _GEN_7; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_9 = 7'h9 == io_ar_addr ? bht_9 : _GEN_8; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_10 = 7'ha == io_ar_addr ? bht_10 : _GEN_9; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_11 = 7'hb == io_ar_addr ? bht_11 : _GEN_10; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_12 = 7'hc == io_ar_addr ? bht_12 : _GEN_11; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_13 = 7'hd == io_ar_addr ? bht_13 : _GEN_12; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_14 = 7'he == io_ar_addr ? bht_14 : _GEN_13; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_15 = 7'hf == io_ar_addr ? bht_15 : _GEN_14; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_16 = 7'h10 == io_ar_addr ? bht_16 : _GEN_15; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_17 = 7'h11 == io_ar_addr ? bht_17 : _GEN_16; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_18 = 7'h12 == io_ar_addr ? bht_18 : _GEN_17; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_19 = 7'h13 == io_ar_addr ? bht_19 : _GEN_18; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_20 = 7'h14 == io_ar_addr ? bht_20 : _GEN_19; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_21 = 7'h15 == io_ar_addr ? bht_21 : _GEN_20; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_22 = 7'h16 == io_ar_addr ? bht_22 : _GEN_21; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_23 = 7'h17 == io_ar_addr ? bht_23 : _GEN_22; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_24 = 7'h18 == io_ar_addr ? bht_24 : _GEN_23; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_25 = 7'h19 == io_ar_addr ? bht_25 : _GEN_24; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_26 = 7'h1a == io_ar_addr ? bht_26 : _GEN_25; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_27 = 7'h1b == io_ar_addr ? bht_27 : _GEN_26; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_28 = 7'h1c == io_ar_addr ? bht_28 : _GEN_27; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_29 = 7'h1d == io_ar_addr ? bht_29 : _GEN_28; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_30 = 7'h1e == io_ar_addr ? bht_30 : _GEN_29; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_31 = 7'h1f == io_ar_addr ? bht_31 : _GEN_30; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_32 = 7'h20 == io_ar_addr ? bht_32 : _GEN_31; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_33 = 7'h21 == io_ar_addr ? bht_33 : _GEN_32; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_34 = 7'h22 == io_ar_addr ? bht_34 : _GEN_33; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_35 = 7'h23 == io_ar_addr ? bht_35 : _GEN_34; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_36 = 7'h24 == io_ar_addr ? bht_36 : _GEN_35; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_37 = 7'h25 == io_ar_addr ? bht_37 : _GEN_36; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_38 = 7'h26 == io_ar_addr ? bht_38 : _GEN_37; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_39 = 7'h27 == io_ar_addr ? bht_39 : _GEN_38; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_40 = 7'h28 == io_ar_addr ? bht_40 : _GEN_39; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_41 = 7'h29 == io_ar_addr ? bht_41 : _GEN_40; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_42 = 7'h2a == io_ar_addr ? bht_42 : _GEN_41; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_43 = 7'h2b == io_ar_addr ? bht_43 : _GEN_42; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_44 = 7'h2c == io_ar_addr ? bht_44 : _GEN_43; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_45 = 7'h2d == io_ar_addr ? bht_45 : _GEN_44; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_46 = 7'h2e == io_ar_addr ? bht_46 : _GEN_45; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_47 = 7'h2f == io_ar_addr ? bht_47 : _GEN_46; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_48 = 7'h30 == io_ar_addr ? bht_48 : _GEN_47; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_49 = 7'h31 == io_ar_addr ? bht_49 : _GEN_48; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_50 = 7'h32 == io_ar_addr ? bht_50 : _GEN_49; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_51 = 7'h33 == io_ar_addr ? bht_51 : _GEN_50; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_52 = 7'h34 == io_ar_addr ? bht_52 : _GEN_51; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_53 = 7'h35 == io_ar_addr ? bht_53 : _GEN_52; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_54 = 7'h36 == io_ar_addr ? bht_54 : _GEN_53; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_55 = 7'h37 == io_ar_addr ? bht_55 : _GEN_54; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_56 = 7'h38 == io_ar_addr ? bht_56 : _GEN_55; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_57 = 7'h39 == io_ar_addr ? bht_57 : _GEN_56; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_58 = 7'h3a == io_ar_addr ? bht_58 : _GEN_57; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_59 = 7'h3b == io_ar_addr ? bht_59 : _GEN_58; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_60 = 7'h3c == io_ar_addr ? bht_60 : _GEN_59; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_61 = 7'h3d == io_ar_addr ? bht_61 : _GEN_60; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_62 = 7'h3e == io_ar_addr ? bht_62 : _GEN_61; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_63 = 7'h3f == io_ar_addr ? bht_63 : _GEN_62; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_64 = 7'h40 == io_ar_addr ? bht_64 : _GEN_63; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_65 = 7'h41 == io_ar_addr ? bht_65 : _GEN_64; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_66 = 7'h42 == io_ar_addr ? bht_66 : _GEN_65; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_67 = 7'h43 == io_ar_addr ? bht_67 : _GEN_66; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_68 = 7'h44 == io_ar_addr ? bht_68 : _GEN_67; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_69 = 7'h45 == io_ar_addr ? bht_69 : _GEN_68; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_70 = 7'h46 == io_ar_addr ? bht_70 : _GEN_69; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_71 = 7'h47 == io_ar_addr ? bht_71 : _GEN_70; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_72 = 7'h48 == io_ar_addr ? bht_72 : _GEN_71; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_73 = 7'h49 == io_ar_addr ? bht_73 : _GEN_72; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_74 = 7'h4a == io_ar_addr ? bht_74 : _GEN_73; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_75 = 7'h4b == io_ar_addr ? bht_75 : _GEN_74; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_76 = 7'h4c == io_ar_addr ? bht_76 : _GEN_75; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_77 = 7'h4d == io_ar_addr ? bht_77 : _GEN_76; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_78 = 7'h4e == io_ar_addr ? bht_78 : _GEN_77; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_79 = 7'h4f == io_ar_addr ? bht_79 : _GEN_78; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_80 = 7'h50 == io_ar_addr ? bht_80 : _GEN_79; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_81 = 7'h51 == io_ar_addr ? bht_81 : _GEN_80; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_82 = 7'h52 == io_ar_addr ? bht_82 : _GEN_81; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_83 = 7'h53 == io_ar_addr ? bht_83 : _GEN_82; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_84 = 7'h54 == io_ar_addr ? bht_84 : _GEN_83; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_85 = 7'h55 == io_ar_addr ? bht_85 : _GEN_84; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_86 = 7'h56 == io_ar_addr ? bht_86 : _GEN_85; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_87 = 7'h57 == io_ar_addr ? bht_87 : _GEN_86; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_88 = 7'h58 == io_ar_addr ? bht_88 : _GEN_87; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_89 = 7'h59 == io_ar_addr ? bht_89 : _GEN_88; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_90 = 7'h5a == io_ar_addr ? bht_90 : _GEN_89; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_91 = 7'h5b == io_ar_addr ? bht_91 : _GEN_90; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_92 = 7'h5c == io_ar_addr ? bht_92 : _GEN_91; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_93 = 7'h5d == io_ar_addr ? bht_93 : _GEN_92; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_94 = 7'h5e == io_ar_addr ? bht_94 : _GEN_93; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_95 = 7'h5f == io_ar_addr ? bht_95 : _GEN_94; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_96 = 7'h60 == io_ar_addr ? bht_96 : _GEN_95; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_97 = 7'h61 == io_ar_addr ? bht_97 : _GEN_96; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_98 = 7'h62 == io_ar_addr ? bht_98 : _GEN_97; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_99 = 7'h63 == io_ar_addr ? bht_99 : _GEN_98; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_100 = 7'h64 == io_ar_addr ? bht_100 : _GEN_99; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_101 = 7'h65 == io_ar_addr ? bht_101 : _GEN_100; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_102 = 7'h66 == io_ar_addr ? bht_102 : _GEN_101; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_103 = 7'h67 == io_ar_addr ? bht_103 : _GEN_102; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_104 = 7'h68 == io_ar_addr ? bht_104 : _GEN_103; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_105 = 7'h69 == io_ar_addr ? bht_105 : _GEN_104; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_106 = 7'h6a == io_ar_addr ? bht_106 : _GEN_105; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_107 = 7'h6b == io_ar_addr ? bht_107 : _GEN_106; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_108 = 7'h6c == io_ar_addr ? bht_108 : _GEN_107; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_109 = 7'h6d == io_ar_addr ? bht_109 : _GEN_108; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_110 = 7'h6e == io_ar_addr ? bht_110 : _GEN_109; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_111 = 7'h6f == io_ar_addr ? bht_111 : _GEN_110; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_112 = 7'h70 == io_ar_addr ? bht_112 : _GEN_111; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_113 = 7'h71 == io_ar_addr ? bht_113 : _GEN_112; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_114 = 7'h72 == io_ar_addr ? bht_114 : _GEN_113; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_115 = 7'h73 == io_ar_addr ? bht_115 : _GEN_114; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_116 = 7'h74 == io_ar_addr ? bht_116 : _GEN_115; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_117 = 7'h75 == io_ar_addr ? bht_117 : _GEN_116; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_118 = 7'h76 == io_ar_addr ? bht_118 : _GEN_117; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_119 = 7'h77 == io_ar_addr ? bht_119 : _GEN_118; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_120 = 7'h78 == io_ar_addr ? bht_120 : _GEN_119; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_121 = 7'h79 == io_ar_addr ? bht_121 : _GEN_120; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_122 = 7'h7a == io_ar_addr ? bht_122 : _GEN_121; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_123 = 7'h7b == io_ar_addr ? bht_123 : _GEN_122; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_124 = 7'h7c == io_ar_addr ? bht_124 : _GEN_123; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_125 = 7'h7d == io_ar_addr ? bht_125 : _GEN_124; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_126 = 7'h7e == io_ar_addr ? bht_126 : _GEN_125; // @[BHT.scala 21:{12,12}]
  assign io_out = 7'h7f == io_ar_addr ? bht_127 : _GEN_126; // @[BHT.scala 21:{12,12}]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_0 <= 3'h0;
    end else if (io_write & 7'h0 == io_aw_addr) begin
      bht_0 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_1 <= 3'h0;
    end else if (io_write & 7'h1 == io_aw_addr) begin
      bht_1 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_2 <= 3'h0;
    end else if (io_write & 7'h2 == io_aw_addr) begin
      bht_2 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_3 <= 3'h0;
    end else if (io_write & 7'h3 == io_aw_addr) begin
      bht_3 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_4 <= 3'h0;
    end else if (io_write & 7'h4 == io_aw_addr) begin
      bht_4 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_5 <= 3'h0;
    end else if (io_write & 7'h5 == io_aw_addr) begin
      bht_5 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_6 <= 3'h0;
    end else if (io_write & 7'h6 == io_aw_addr) begin
      bht_6 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_7 <= 3'h0;
    end else if (io_write & 7'h7 == io_aw_addr) begin
      bht_7 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_8 <= 3'h0;
    end else if (io_write & 7'h8 == io_aw_addr) begin
      bht_8 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_9 <= 3'h0;
    end else if (io_write & 7'h9 == io_aw_addr) begin
      bht_9 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_10 <= 3'h0;
    end else if (io_write & 7'ha == io_aw_addr) begin
      bht_10 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_11 <= 3'h0;
    end else if (io_write & 7'hb == io_aw_addr) begin
      bht_11 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_12 <= 3'h0;
    end else if (io_write & 7'hc == io_aw_addr) begin
      bht_12 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_13 <= 3'h0;
    end else if (io_write & 7'hd == io_aw_addr) begin
      bht_13 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_14 <= 3'h0;
    end else if (io_write & 7'he == io_aw_addr) begin
      bht_14 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_15 <= 3'h0;
    end else if (io_write & 7'hf == io_aw_addr) begin
      bht_15 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_16 <= 3'h0;
    end else if (io_write & 7'h10 == io_aw_addr) begin
      bht_16 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_17 <= 3'h0;
    end else if (io_write & 7'h11 == io_aw_addr) begin
      bht_17 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_18 <= 3'h0;
    end else if (io_write & 7'h12 == io_aw_addr) begin
      bht_18 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_19 <= 3'h0;
    end else if (io_write & 7'h13 == io_aw_addr) begin
      bht_19 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_20 <= 3'h0;
    end else if (io_write & 7'h14 == io_aw_addr) begin
      bht_20 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_21 <= 3'h0;
    end else if (io_write & 7'h15 == io_aw_addr) begin
      bht_21 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_22 <= 3'h0;
    end else if (io_write & 7'h16 == io_aw_addr) begin
      bht_22 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_23 <= 3'h0;
    end else if (io_write & 7'h17 == io_aw_addr) begin
      bht_23 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_24 <= 3'h0;
    end else if (io_write & 7'h18 == io_aw_addr) begin
      bht_24 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_25 <= 3'h0;
    end else if (io_write & 7'h19 == io_aw_addr) begin
      bht_25 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_26 <= 3'h0;
    end else if (io_write & 7'h1a == io_aw_addr) begin
      bht_26 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_27 <= 3'h0;
    end else if (io_write & 7'h1b == io_aw_addr) begin
      bht_27 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_28 <= 3'h0;
    end else if (io_write & 7'h1c == io_aw_addr) begin
      bht_28 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_29 <= 3'h0;
    end else if (io_write & 7'h1d == io_aw_addr) begin
      bht_29 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_30 <= 3'h0;
    end else if (io_write & 7'h1e == io_aw_addr) begin
      bht_30 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_31 <= 3'h0;
    end else if (io_write & 7'h1f == io_aw_addr) begin
      bht_31 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_32 <= 3'h0;
    end else if (io_write & 7'h20 == io_aw_addr) begin
      bht_32 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_33 <= 3'h0;
    end else if (io_write & 7'h21 == io_aw_addr) begin
      bht_33 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_34 <= 3'h0;
    end else if (io_write & 7'h22 == io_aw_addr) begin
      bht_34 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_35 <= 3'h0;
    end else if (io_write & 7'h23 == io_aw_addr) begin
      bht_35 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_36 <= 3'h0;
    end else if (io_write & 7'h24 == io_aw_addr) begin
      bht_36 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_37 <= 3'h0;
    end else if (io_write & 7'h25 == io_aw_addr) begin
      bht_37 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_38 <= 3'h0;
    end else if (io_write & 7'h26 == io_aw_addr) begin
      bht_38 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_39 <= 3'h0;
    end else if (io_write & 7'h27 == io_aw_addr) begin
      bht_39 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_40 <= 3'h0;
    end else if (io_write & 7'h28 == io_aw_addr) begin
      bht_40 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_41 <= 3'h0;
    end else if (io_write & 7'h29 == io_aw_addr) begin
      bht_41 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_42 <= 3'h0;
    end else if (io_write & 7'h2a == io_aw_addr) begin
      bht_42 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_43 <= 3'h0;
    end else if (io_write & 7'h2b == io_aw_addr) begin
      bht_43 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_44 <= 3'h0;
    end else if (io_write & 7'h2c == io_aw_addr) begin
      bht_44 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_45 <= 3'h0;
    end else if (io_write & 7'h2d == io_aw_addr) begin
      bht_45 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_46 <= 3'h0;
    end else if (io_write & 7'h2e == io_aw_addr) begin
      bht_46 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_47 <= 3'h0;
    end else if (io_write & 7'h2f == io_aw_addr) begin
      bht_47 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_48 <= 3'h0;
    end else if (io_write & 7'h30 == io_aw_addr) begin
      bht_48 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_49 <= 3'h0;
    end else if (io_write & 7'h31 == io_aw_addr) begin
      bht_49 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_50 <= 3'h0;
    end else if (io_write & 7'h32 == io_aw_addr) begin
      bht_50 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_51 <= 3'h0;
    end else if (io_write & 7'h33 == io_aw_addr) begin
      bht_51 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_52 <= 3'h0;
    end else if (io_write & 7'h34 == io_aw_addr) begin
      bht_52 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_53 <= 3'h0;
    end else if (io_write & 7'h35 == io_aw_addr) begin
      bht_53 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_54 <= 3'h0;
    end else if (io_write & 7'h36 == io_aw_addr) begin
      bht_54 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_55 <= 3'h0;
    end else if (io_write & 7'h37 == io_aw_addr) begin
      bht_55 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_56 <= 3'h0;
    end else if (io_write & 7'h38 == io_aw_addr) begin
      bht_56 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_57 <= 3'h0;
    end else if (io_write & 7'h39 == io_aw_addr) begin
      bht_57 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_58 <= 3'h0;
    end else if (io_write & 7'h3a == io_aw_addr) begin
      bht_58 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_59 <= 3'h0;
    end else if (io_write & 7'h3b == io_aw_addr) begin
      bht_59 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_60 <= 3'h0;
    end else if (io_write & 7'h3c == io_aw_addr) begin
      bht_60 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_61 <= 3'h0;
    end else if (io_write & 7'h3d == io_aw_addr) begin
      bht_61 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_62 <= 3'h0;
    end else if (io_write & 7'h3e == io_aw_addr) begin
      bht_62 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_63 <= 3'h0;
    end else if (io_write & 7'h3f == io_aw_addr) begin
      bht_63 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_64 <= 3'h0;
    end else if (io_write & 7'h40 == io_aw_addr) begin
      bht_64 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_65 <= 3'h0;
    end else if (io_write & 7'h41 == io_aw_addr) begin
      bht_65 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_66 <= 3'h0;
    end else if (io_write & 7'h42 == io_aw_addr) begin
      bht_66 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_67 <= 3'h0;
    end else if (io_write & 7'h43 == io_aw_addr) begin
      bht_67 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_68 <= 3'h0;
    end else if (io_write & 7'h44 == io_aw_addr) begin
      bht_68 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_69 <= 3'h0;
    end else if (io_write & 7'h45 == io_aw_addr) begin
      bht_69 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_70 <= 3'h0;
    end else if (io_write & 7'h46 == io_aw_addr) begin
      bht_70 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_71 <= 3'h0;
    end else if (io_write & 7'h47 == io_aw_addr) begin
      bht_71 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_72 <= 3'h0;
    end else if (io_write & 7'h48 == io_aw_addr) begin
      bht_72 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_73 <= 3'h0;
    end else if (io_write & 7'h49 == io_aw_addr) begin
      bht_73 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_74 <= 3'h0;
    end else if (io_write & 7'h4a == io_aw_addr) begin
      bht_74 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_75 <= 3'h0;
    end else if (io_write & 7'h4b == io_aw_addr) begin
      bht_75 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_76 <= 3'h0;
    end else if (io_write & 7'h4c == io_aw_addr) begin
      bht_76 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_77 <= 3'h0;
    end else if (io_write & 7'h4d == io_aw_addr) begin
      bht_77 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_78 <= 3'h0;
    end else if (io_write & 7'h4e == io_aw_addr) begin
      bht_78 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_79 <= 3'h0;
    end else if (io_write & 7'h4f == io_aw_addr) begin
      bht_79 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_80 <= 3'h0;
    end else if (io_write & 7'h50 == io_aw_addr) begin
      bht_80 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_81 <= 3'h0;
    end else if (io_write & 7'h51 == io_aw_addr) begin
      bht_81 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_82 <= 3'h0;
    end else if (io_write & 7'h52 == io_aw_addr) begin
      bht_82 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_83 <= 3'h0;
    end else if (io_write & 7'h53 == io_aw_addr) begin
      bht_83 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_84 <= 3'h0;
    end else if (io_write & 7'h54 == io_aw_addr) begin
      bht_84 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_85 <= 3'h0;
    end else if (io_write & 7'h55 == io_aw_addr) begin
      bht_85 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_86 <= 3'h0;
    end else if (io_write & 7'h56 == io_aw_addr) begin
      bht_86 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_87 <= 3'h0;
    end else if (io_write & 7'h57 == io_aw_addr) begin
      bht_87 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_88 <= 3'h0;
    end else if (io_write & 7'h58 == io_aw_addr) begin
      bht_88 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_89 <= 3'h0;
    end else if (io_write & 7'h59 == io_aw_addr) begin
      bht_89 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_90 <= 3'h0;
    end else if (io_write & 7'h5a == io_aw_addr) begin
      bht_90 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_91 <= 3'h0;
    end else if (io_write & 7'h5b == io_aw_addr) begin
      bht_91 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_92 <= 3'h0;
    end else if (io_write & 7'h5c == io_aw_addr) begin
      bht_92 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_93 <= 3'h0;
    end else if (io_write & 7'h5d == io_aw_addr) begin
      bht_93 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_94 <= 3'h0;
    end else if (io_write & 7'h5e == io_aw_addr) begin
      bht_94 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_95 <= 3'h0;
    end else if (io_write & 7'h5f == io_aw_addr) begin
      bht_95 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_96 <= 3'h0;
    end else if (io_write & 7'h60 == io_aw_addr) begin
      bht_96 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_97 <= 3'h0;
    end else if (io_write & 7'h61 == io_aw_addr) begin
      bht_97 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_98 <= 3'h0;
    end else if (io_write & 7'h62 == io_aw_addr) begin
      bht_98 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_99 <= 3'h0;
    end else if (io_write & 7'h63 == io_aw_addr) begin
      bht_99 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_100 <= 3'h0;
    end else if (io_write & 7'h64 == io_aw_addr) begin
      bht_100 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_101 <= 3'h0;
    end else if (io_write & 7'h65 == io_aw_addr) begin
      bht_101 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_102 <= 3'h0;
    end else if (io_write & 7'h66 == io_aw_addr) begin
      bht_102 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_103 <= 3'h0;
    end else if (io_write & 7'h67 == io_aw_addr) begin
      bht_103 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_104 <= 3'h0;
    end else if (io_write & 7'h68 == io_aw_addr) begin
      bht_104 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_105 <= 3'h0;
    end else if (io_write & 7'h69 == io_aw_addr) begin
      bht_105 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_106 <= 3'h0;
    end else if (io_write & 7'h6a == io_aw_addr) begin
      bht_106 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_107 <= 3'h0;
    end else if (io_write & 7'h6b == io_aw_addr) begin
      bht_107 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_108 <= 3'h0;
    end else if (io_write & 7'h6c == io_aw_addr) begin
      bht_108 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_109 <= 3'h0;
    end else if (io_write & 7'h6d == io_aw_addr) begin
      bht_109 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_110 <= 3'h0;
    end else if (io_write & 7'h6e == io_aw_addr) begin
      bht_110 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_111 <= 3'h0;
    end else if (io_write & 7'h6f == io_aw_addr) begin
      bht_111 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_112 <= 3'h0;
    end else if (io_write & 7'h70 == io_aw_addr) begin
      bht_112 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_113 <= 3'h0;
    end else if (io_write & 7'h71 == io_aw_addr) begin
      bht_113 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_114 <= 3'h0;
    end else if (io_write & 7'h72 == io_aw_addr) begin
      bht_114 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_115 <= 3'h0;
    end else if (io_write & 7'h73 == io_aw_addr) begin
      bht_115 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_116 <= 3'h0;
    end else if (io_write & 7'h74 == io_aw_addr) begin
      bht_116 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_117 <= 3'h0;
    end else if (io_write & 7'h75 == io_aw_addr) begin
      bht_117 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_118 <= 3'h0;
    end else if (io_write & 7'h76 == io_aw_addr) begin
      bht_118 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_119 <= 3'h0;
    end else if (io_write & 7'h77 == io_aw_addr) begin
      bht_119 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_120 <= 3'h0;
    end else if (io_write & 7'h78 == io_aw_addr) begin
      bht_120 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_121 <= 3'h0;
    end else if (io_write & 7'h79 == io_aw_addr) begin
      bht_121 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_122 <= 3'h0;
    end else if (io_write & 7'h7a == io_aw_addr) begin
      bht_122 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_123 <= 3'h0;
    end else if (io_write & 7'h7b == io_aw_addr) begin
      bht_123 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_124 <= 3'h0;
    end else if (io_write & 7'h7c == io_aw_addr) begin
      bht_124 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_125 <= 3'h0;
    end else if (io_write & 7'h7d == io_aw_addr) begin
      bht_125 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_126 <= 3'h0;
    end else if (io_write & 7'h7e == io_aw_addr) begin
      bht_126 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_127 <= 3'h0;
    end else if (io_write & 7'h7f == io_aw_addr) begin
      bht_127 <= io_in;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bht_0 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bht_1 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  bht_2 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  bht_3 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  bht_4 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  bht_5 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  bht_6 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  bht_7 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  bht_8 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  bht_9 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  bht_10 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  bht_11 = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  bht_12 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  bht_13 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  bht_14 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  bht_15 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  bht_16 = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  bht_17 = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  bht_18 = _RAND_18[2:0];
  _RAND_19 = {1{`RANDOM}};
  bht_19 = _RAND_19[2:0];
  _RAND_20 = {1{`RANDOM}};
  bht_20 = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  bht_21 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  bht_22 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  bht_23 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  bht_24 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  bht_25 = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  bht_26 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  bht_27 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  bht_28 = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  bht_29 = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  bht_30 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  bht_31 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  bht_32 = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  bht_33 = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  bht_34 = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  bht_35 = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  bht_36 = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  bht_37 = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  bht_38 = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  bht_39 = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  bht_40 = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  bht_41 = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  bht_42 = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  bht_43 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  bht_44 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  bht_45 = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  bht_46 = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  bht_47 = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  bht_48 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  bht_49 = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  bht_50 = _RAND_50[2:0];
  _RAND_51 = {1{`RANDOM}};
  bht_51 = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  bht_52 = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  bht_53 = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  bht_54 = _RAND_54[2:0];
  _RAND_55 = {1{`RANDOM}};
  bht_55 = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  bht_56 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  bht_57 = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  bht_58 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  bht_59 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  bht_60 = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  bht_61 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  bht_62 = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  bht_63 = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  bht_64 = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  bht_65 = _RAND_65[2:0];
  _RAND_66 = {1{`RANDOM}};
  bht_66 = _RAND_66[2:0];
  _RAND_67 = {1{`RANDOM}};
  bht_67 = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  bht_68 = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  bht_69 = _RAND_69[2:0];
  _RAND_70 = {1{`RANDOM}};
  bht_70 = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  bht_71 = _RAND_71[2:0];
  _RAND_72 = {1{`RANDOM}};
  bht_72 = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  bht_73 = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  bht_74 = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  bht_75 = _RAND_75[2:0];
  _RAND_76 = {1{`RANDOM}};
  bht_76 = _RAND_76[2:0];
  _RAND_77 = {1{`RANDOM}};
  bht_77 = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  bht_78 = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  bht_79 = _RAND_79[2:0];
  _RAND_80 = {1{`RANDOM}};
  bht_80 = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  bht_81 = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  bht_82 = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  bht_83 = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  bht_84 = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  bht_85 = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  bht_86 = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  bht_87 = _RAND_87[2:0];
  _RAND_88 = {1{`RANDOM}};
  bht_88 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  bht_89 = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  bht_90 = _RAND_90[2:0];
  _RAND_91 = {1{`RANDOM}};
  bht_91 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  bht_92 = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  bht_93 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  bht_94 = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  bht_95 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  bht_96 = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  bht_97 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  bht_98 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  bht_99 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  bht_100 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  bht_101 = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  bht_102 = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  bht_103 = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  bht_104 = _RAND_104[2:0];
  _RAND_105 = {1{`RANDOM}};
  bht_105 = _RAND_105[2:0];
  _RAND_106 = {1{`RANDOM}};
  bht_106 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  bht_107 = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  bht_108 = _RAND_108[2:0];
  _RAND_109 = {1{`RANDOM}};
  bht_109 = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  bht_110 = _RAND_110[2:0];
  _RAND_111 = {1{`RANDOM}};
  bht_111 = _RAND_111[2:0];
  _RAND_112 = {1{`RANDOM}};
  bht_112 = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  bht_113 = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  bht_114 = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  bht_115 = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  bht_116 = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  bht_117 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  bht_118 = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  bht_119 = _RAND_119[2:0];
  _RAND_120 = {1{`RANDOM}};
  bht_120 = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  bht_121 = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  bht_122 = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  bht_123 = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  bht_124 = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  bht_125 = _RAND_125[2:0];
  _RAND_126 = {1{`RANDOM}};
  bht_126 = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  bht_127 = _RAND_127[2:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    bht_0 = 3'h0;
  end
  if (reset) begin
    bht_1 = 3'h0;
  end
  if (reset) begin
    bht_2 = 3'h0;
  end
  if (reset) begin
    bht_3 = 3'h0;
  end
  if (reset) begin
    bht_4 = 3'h0;
  end
  if (reset) begin
    bht_5 = 3'h0;
  end
  if (reset) begin
    bht_6 = 3'h0;
  end
  if (reset) begin
    bht_7 = 3'h0;
  end
  if (reset) begin
    bht_8 = 3'h0;
  end
  if (reset) begin
    bht_9 = 3'h0;
  end
  if (reset) begin
    bht_10 = 3'h0;
  end
  if (reset) begin
    bht_11 = 3'h0;
  end
  if (reset) begin
    bht_12 = 3'h0;
  end
  if (reset) begin
    bht_13 = 3'h0;
  end
  if (reset) begin
    bht_14 = 3'h0;
  end
  if (reset) begin
    bht_15 = 3'h0;
  end
  if (reset) begin
    bht_16 = 3'h0;
  end
  if (reset) begin
    bht_17 = 3'h0;
  end
  if (reset) begin
    bht_18 = 3'h0;
  end
  if (reset) begin
    bht_19 = 3'h0;
  end
  if (reset) begin
    bht_20 = 3'h0;
  end
  if (reset) begin
    bht_21 = 3'h0;
  end
  if (reset) begin
    bht_22 = 3'h0;
  end
  if (reset) begin
    bht_23 = 3'h0;
  end
  if (reset) begin
    bht_24 = 3'h0;
  end
  if (reset) begin
    bht_25 = 3'h0;
  end
  if (reset) begin
    bht_26 = 3'h0;
  end
  if (reset) begin
    bht_27 = 3'h0;
  end
  if (reset) begin
    bht_28 = 3'h0;
  end
  if (reset) begin
    bht_29 = 3'h0;
  end
  if (reset) begin
    bht_30 = 3'h0;
  end
  if (reset) begin
    bht_31 = 3'h0;
  end
  if (reset) begin
    bht_32 = 3'h0;
  end
  if (reset) begin
    bht_33 = 3'h0;
  end
  if (reset) begin
    bht_34 = 3'h0;
  end
  if (reset) begin
    bht_35 = 3'h0;
  end
  if (reset) begin
    bht_36 = 3'h0;
  end
  if (reset) begin
    bht_37 = 3'h0;
  end
  if (reset) begin
    bht_38 = 3'h0;
  end
  if (reset) begin
    bht_39 = 3'h0;
  end
  if (reset) begin
    bht_40 = 3'h0;
  end
  if (reset) begin
    bht_41 = 3'h0;
  end
  if (reset) begin
    bht_42 = 3'h0;
  end
  if (reset) begin
    bht_43 = 3'h0;
  end
  if (reset) begin
    bht_44 = 3'h0;
  end
  if (reset) begin
    bht_45 = 3'h0;
  end
  if (reset) begin
    bht_46 = 3'h0;
  end
  if (reset) begin
    bht_47 = 3'h0;
  end
  if (reset) begin
    bht_48 = 3'h0;
  end
  if (reset) begin
    bht_49 = 3'h0;
  end
  if (reset) begin
    bht_50 = 3'h0;
  end
  if (reset) begin
    bht_51 = 3'h0;
  end
  if (reset) begin
    bht_52 = 3'h0;
  end
  if (reset) begin
    bht_53 = 3'h0;
  end
  if (reset) begin
    bht_54 = 3'h0;
  end
  if (reset) begin
    bht_55 = 3'h0;
  end
  if (reset) begin
    bht_56 = 3'h0;
  end
  if (reset) begin
    bht_57 = 3'h0;
  end
  if (reset) begin
    bht_58 = 3'h0;
  end
  if (reset) begin
    bht_59 = 3'h0;
  end
  if (reset) begin
    bht_60 = 3'h0;
  end
  if (reset) begin
    bht_61 = 3'h0;
  end
  if (reset) begin
    bht_62 = 3'h0;
  end
  if (reset) begin
    bht_63 = 3'h0;
  end
  if (reset) begin
    bht_64 = 3'h0;
  end
  if (reset) begin
    bht_65 = 3'h0;
  end
  if (reset) begin
    bht_66 = 3'h0;
  end
  if (reset) begin
    bht_67 = 3'h0;
  end
  if (reset) begin
    bht_68 = 3'h0;
  end
  if (reset) begin
    bht_69 = 3'h0;
  end
  if (reset) begin
    bht_70 = 3'h0;
  end
  if (reset) begin
    bht_71 = 3'h0;
  end
  if (reset) begin
    bht_72 = 3'h0;
  end
  if (reset) begin
    bht_73 = 3'h0;
  end
  if (reset) begin
    bht_74 = 3'h0;
  end
  if (reset) begin
    bht_75 = 3'h0;
  end
  if (reset) begin
    bht_76 = 3'h0;
  end
  if (reset) begin
    bht_77 = 3'h0;
  end
  if (reset) begin
    bht_78 = 3'h0;
  end
  if (reset) begin
    bht_79 = 3'h0;
  end
  if (reset) begin
    bht_80 = 3'h0;
  end
  if (reset) begin
    bht_81 = 3'h0;
  end
  if (reset) begin
    bht_82 = 3'h0;
  end
  if (reset) begin
    bht_83 = 3'h0;
  end
  if (reset) begin
    bht_84 = 3'h0;
  end
  if (reset) begin
    bht_85 = 3'h0;
  end
  if (reset) begin
    bht_86 = 3'h0;
  end
  if (reset) begin
    bht_87 = 3'h0;
  end
  if (reset) begin
    bht_88 = 3'h0;
  end
  if (reset) begin
    bht_89 = 3'h0;
  end
  if (reset) begin
    bht_90 = 3'h0;
  end
  if (reset) begin
    bht_91 = 3'h0;
  end
  if (reset) begin
    bht_92 = 3'h0;
  end
  if (reset) begin
    bht_93 = 3'h0;
  end
  if (reset) begin
    bht_94 = 3'h0;
  end
  if (reset) begin
    bht_95 = 3'h0;
  end
  if (reset) begin
    bht_96 = 3'h0;
  end
  if (reset) begin
    bht_97 = 3'h0;
  end
  if (reset) begin
    bht_98 = 3'h0;
  end
  if (reset) begin
    bht_99 = 3'h0;
  end
  if (reset) begin
    bht_100 = 3'h0;
  end
  if (reset) begin
    bht_101 = 3'h0;
  end
  if (reset) begin
    bht_102 = 3'h0;
  end
  if (reset) begin
    bht_103 = 3'h0;
  end
  if (reset) begin
    bht_104 = 3'h0;
  end
  if (reset) begin
    bht_105 = 3'h0;
  end
  if (reset) begin
    bht_106 = 3'h0;
  end
  if (reset) begin
    bht_107 = 3'h0;
  end
  if (reset) begin
    bht_108 = 3'h0;
  end
  if (reset) begin
    bht_109 = 3'h0;
  end
  if (reset) begin
    bht_110 = 3'h0;
  end
  if (reset) begin
    bht_111 = 3'h0;
  end
  if (reset) begin
    bht_112 = 3'h0;
  end
  if (reset) begin
    bht_113 = 3'h0;
  end
  if (reset) begin
    bht_114 = 3'h0;
  end
  if (reset) begin
    bht_115 = 3'h0;
  end
  if (reset) begin
    bht_116 = 3'h0;
  end
  if (reset) begin
    bht_117 = 3'h0;
  end
  if (reset) begin
    bht_118 = 3'h0;
  end
  if (reset) begin
    bht_119 = 3'h0;
  end
  if (reset) begin
    bht_120 = 3'h0;
  end
  if (reset) begin
    bht_121 = 3'h0;
  end
  if (reset) begin
    bht_122 = 3'h0;
  end
  if (reset) begin
    bht_123 = 3'h0;
  end
  if (reset) begin
    bht_124 = 3'h0;
  end
  if (reset) begin
    bht_125 = 3'h0;
  end
  if (reset) begin
    bht_126 = 3'h0;
  end
  if (reset) begin
    bht_127 = 3'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BHT_banks_oneissue(
  input        clock,
  input        reset,
  input  [1:0] io_ar_bank_sel,
  input  [6:0] io_ar_addr_L,
  input  [6:0] io_aw_addr,
  input        io_write,
  input  [2:0] io_in,
  output [2:0] io_out_L
);
  wire  BHT_clock; // @[BHT.scala 84:54]
  wire  BHT_reset; // @[BHT.scala 84:54]
  wire [6:0] BHT_io_ar_addr; // @[BHT.scala 84:54]
  wire [6:0] BHT_io_aw_addr; // @[BHT.scala 84:54]
  wire  BHT_io_write; // @[BHT.scala 84:54]
  wire [2:0] BHT_io_in; // @[BHT.scala 84:54]
  wire [2:0] BHT_io_out; // @[BHT.scala 84:54]
  wire  BHT_1_clock; // @[BHT.scala 84:54]
  wire  BHT_1_reset; // @[BHT.scala 84:54]
  wire [6:0] BHT_1_io_ar_addr; // @[BHT.scala 84:54]
  wire [6:0] BHT_1_io_aw_addr; // @[BHT.scala 84:54]
  wire  BHT_1_io_write; // @[BHT.scala 84:54]
  wire [2:0] BHT_1_io_in; // @[BHT.scala 84:54]
  wire [2:0] BHT_1_io_out; // @[BHT.scala 84:54]
  wire  BHT_2_clock; // @[BHT.scala 84:54]
  wire  BHT_2_reset; // @[BHT.scala 84:54]
  wire [6:0] BHT_2_io_ar_addr; // @[BHT.scala 84:54]
  wire [6:0] BHT_2_io_aw_addr; // @[BHT.scala 84:54]
  wire  BHT_2_io_write; // @[BHT.scala 84:54]
  wire [2:0] BHT_2_io_in; // @[BHT.scala 84:54]
  wire [2:0] BHT_2_io_out; // @[BHT.scala 84:54]
  wire  BHT_3_clock; // @[BHT.scala 84:54]
  wire  BHT_3_reset; // @[BHT.scala 84:54]
  wire [6:0] BHT_3_io_ar_addr; // @[BHT.scala 84:54]
  wire [6:0] BHT_3_io_aw_addr; // @[BHT.scala 84:54]
  wire  BHT_3_io_write; // @[BHT.scala 84:54]
  wire [2:0] BHT_3_io_in; // @[BHT.scala 84:54]
  wire [2:0] BHT_3_io_out; // @[BHT.scala 84:54]
  wire [2:0] bht_banks_0_out = BHT_io_out; // @[BHT.scala 84:{28,28}]
  wire [2:0] bht_banks_1_out = BHT_1_io_out; // @[BHT.scala 84:{28,28}]
  wire [2:0] _GEN_1 = 2'h1 == io_ar_bank_sel ? bht_banks_1_out : bht_banks_0_out; // @[BHT.scala 96:{14,14}]
  wire [2:0] bht_banks_2_out = BHT_2_io_out; // @[BHT.scala 84:{28,28}]
  wire [2:0] _GEN_2 = 2'h2 == io_ar_bank_sel ? bht_banks_2_out : _GEN_1; // @[BHT.scala 96:{14,14}]
  wire [2:0] bht_banks_3_out = BHT_3_io_out; // @[BHT.scala 84:{28,28}]
  BHT BHT ( // @[BHT.scala 84:54]
    .clock(BHT_clock),
    .reset(BHT_reset),
    .io_ar_addr(BHT_io_ar_addr),
    .io_aw_addr(BHT_io_aw_addr),
    .io_write(BHT_io_write),
    .io_in(BHT_io_in),
    .io_out(BHT_io_out)
  );
  BHT BHT_1 ( // @[BHT.scala 84:54]
    .clock(BHT_1_clock),
    .reset(BHT_1_reset),
    .io_ar_addr(BHT_1_io_ar_addr),
    .io_aw_addr(BHT_1_io_aw_addr),
    .io_write(BHT_1_io_write),
    .io_in(BHT_1_io_in),
    .io_out(BHT_1_io_out)
  );
  BHT BHT_2 ( // @[BHT.scala 84:54]
    .clock(BHT_2_clock),
    .reset(BHT_2_reset),
    .io_ar_addr(BHT_2_io_ar_addr),
    .io_aw_addr(BHT_2_io_aw_addr),
    .io_write(BHT_2_io_write),
    .io_in(BHT_2_io_in),
    .io_out(BHT_2_io_out)
  );
  BHT BHT_3 ( // @[BHT.scala 84:54]
    .clock(BHT_3_clock),
    .reset(BHT_3_reset),
    .io_ar_addr(BHT_3_io_ar_addr),
    .io_aw_addr(BHT_3_io_aw_addr),
    .io_write(BHT_3_io_write),
    .io_in(BHT_3_io_in),
    .io_out(BHT_3_io_out)
  );
  assign io_out_L = 2'h3 == io_ar_bank_sel ? bht_banks_3_out : _GEN_2; // @[BHT.scala 96:{14,14}]
  assign BHT_clock = clock;
  assign BHT_reset = reset;
  assign BHT_io_ar_addr = io_ar_addr_L; // @[BHT.scala 84:28 88:30]
  assign BHT_io_aw_addr = io_aw_addr; // @[BHT.scala 84:28 94:30]
  assign BHT_io_write = io_ar_bank_sel == 2'h0 & io_write; // @[BHT.scala 86:59]
  assign BHT_io_in = io_in; // @[BHT.scala 84:28 87:25]
  assign BHT_1_clock = clock;
  assign BHT_1_reset = reset;
  assign BHT_1_io_ar_addr = io_ar_addr_L; // @[BHT.scala 84:28 88:30]
  assign BHT_1_io_aw_addr = io_aw_addr; // @[BHT.scala 84:28 94:30]
  assign BHT_1_io_write = io_ar_bank_sel == 2'h1 & io_write; // @[BHT.scala 86:59]
  assign BHT_1_io_in = io_in; // @[BHT.scala 84:28 87:25]
  assign BHT_2_clock = clock;
  assign BHT_2_reset = reset;
  assign BHT_2_io_ar_addr = io_ar_addr_L; // @[BHT.scala 84:28 88:30]
  assign BHT_2_io_aw_addr = io_aw_addr; // @[BHT.scala 84:28 94:30]
  assign BHT_2_io_write = io_ar_bank_sel == 2'h2 & io_write; // @[BHT.scala 86:59]
  assign BHT_2_io_in = io_in; // @[BHT.scala 84:28 87:25]
  assign BHT_3_clock = clock;
  assign BHT_3_reset = reset;
  assign BHT_3_io_ar_addr = io_ar_addr_L; // @[BHT.scala 84:28 88:30]
  assign BHT_3_io_aw_addr = io_aw_addr; // @[BHT.scala 84:28 94:30]
  assign BHT_3_io_write = io_ar_bank_sel == 2'h3 & io_write; // @[BHT.scala 86:59]
  assign BHT_3_io_in = io_in; // @[BHT.scala 84:28 87:25]
endmodule
module btb_tag_with_block_ram(
  input        clock,
  input        io_wen,
  input  [8:0] io_raddr,
  input  [8:0] io_waddr,
  input  [7:0] io_wdata,
  output [7:0] io_rdata
);
  wire  btb_tag_ram_0_clka; // @[BTB.scala 216:31]
  wire  btb_tag_ram_0_clkb; // @[BTB.scala 216:31]
  wire  btb_tag_ram_0_ena; // @[BTB.scala 216:31]
  wire  btb_tag_ram_0_enb; // @[BTB.scala 216:31]
  wire  btb_tag_ram_0_wea; // @[BTB.scala 216:31]
  wire [8:0] btb_tag_ram_0_addra; // @[BTB.scala 216:31]
  wire [7:0] btb_tag_ram_0_dina; // @[BTB.scala 216:31]
  wire [8:0] btb_tag_ram_0_addrb; // @[BTB.scala 216:31]
  wire [7:0] btb_tag_ram_0_doutb; // @[BTB.scala 216:31]
  btb_tag_ram btb_tag_ram_0 ( // @[BTB.scala 216:31]
    .clka(btb_tag_ram_0_clka),
    .clkb(btb_tag_ram_0_clkb),
    .ena(btb_tag_ram_0_ena),
    .enb(btb_tag_ram_0_enb),
    .wea(btb_tag_ram_0_wea),
    .addra(btb_tag_ram_0_addra),
    .dina(btb_tag_ram_0_dina),
    .addrb(btb_tag_ram_0_addrb),
    .doutb(btb_tag_ram_0_doutb)
  );
  assign io_rdata = btb_tag_ram_0_doutb; // @[BTB.scala 225:18]
  assign btb_tag_ram_0_clka = clock; // @[BTB.scala 217:36]
  assign btb_tag_ram_0_clkb = clock; // @[BTB.scala 218:36]
  assign btb_tag_ram_0_ena = 1'h1; // @[BTB.scala 219:28]
  assign btb_tag_ram_0_enb = 1'h1; // @[BTB.scala 220:28]
  assign btb_tag_ram_0_wea = io_wen; // @[BTB.scala 221:27]
  assign btb_tag_ram_0_addra = io_waddr; // @[BTB.scala 222:28]
  assign btb_tag_ram_0_dina = io_wdata; // @[BTB.scala 224:27]
  assign btb_tag_ram_0_addrb = io_raddr; // @[BTB.scala 223:28]
endmodule
module btb_data_with_block_ram(
  input         clock,
  input         io_wen,
  input  [8:0]  io_raddr,
  input  [8:0]  io_waddr,
  input  [31:0] io_wdata,
  output [31:0] io_rdata
);
  wire  btb_data_ram_0_clka; // @[BTB.scala 189:32]
  wire  btb_data_ram_0_clkb; // @[BTB.scala 189:32]
  wire  btb_data_ram_0_ena; // @[BTB.scala 189:32]
  wire  btb_data_ram_0_enb; // @[BTB.scala 189:32]
  wire  btb_data_ram_0_wea; // @[BTB.scala 189:32]
  wire [8:0] btb_data_ram_0_addra; // @[BTB.scala 189:32]
  wire [31:0] btb_data_ram_0_dina; // @[BTB.scala 189:32]
  wire [8:0] btb_data_ram_0_addrb; // @[BTB.scala 189:32]
  wire [31:0] btb_data_ram_0_doutb; // @[BTB.scala 189:32]
  btb_data_ram btb_data_ram_0 ( // @[BTB.scala 189:32]
    .clka(btb_data_ram_0_clka),
    .clkb(btb_data_ram_0_clkb),
    .ena(btb_data_ram_0_ena),
    .enb(btb_data_ram_0_enb),
    .wea(btb_data_ram_0_wea),
    .addra(btb_data_ram_0_addra),
    .dina(btb_data_ram_0_dina),
    .addrb(btb_data_ram_0_addrb),
    .doutb(btb_data_ram_0_doutb)
  );
  assign io_rdata = btb_data_ram_0_doutb; // @[BTB.scala 198:18]
  assign btb_data_ram_0_clka = clock; // @[BTB.scala 190:37]
  assign btb_data_ram_0_clkb = clock; // @[BTB.scala 191:37]
  assign btb_data_ram_0_ena = 1'h1; // @[BTB.scala 192:29]
  assign btb_data_ram_0_enb = 1'h1; // @[BTB.scala 193:29]
  assign btb_data_ram_0_wea = io_wen; // @[BTB.scala 194:28]
  assign btb_data_ram_0_addra = io_waddr; // @[BTB.scala 195:29]
  assign btb_data_ram_0_dina = io_wdata; // @[BTB.scala 197:28]
  assign btb_data_ram_0_addrb = io_raddr; // @[BTB.scala 196:29]
endmodule
module BTB_banks_oneissue_with_block_ram(
  input         clock,
  input         reset,
  input  [31:0] io_ar_addr_L,
  input  [31:0] io_aw_addr,
  input  [31:0] io_aw_target_addr,
  input         io_write,
  output [31:0] io_out_L,
  output        io_hit_L
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  btb_tag_with_block_ram_clock; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_io_wen; // @[BTB.scala 249:54]
  wire [8:0] btb_tag_with_block_ram_io_raddr; // @[BTB.scala 249:54]
  wire [8:0] btb_tag_with_block_ram_io_waddr; // @[BTB.scala 249:54]
  wire [7:0] btb_tag_with_block_ram_io_wdata; // @[BTB.scala 249:54]
  wire [7:0] btb_tag_with_block_ram_io_rdata; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_1_clock; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_1_io_wen; // @[BTB.scala 249:54]
  wire [8:0] btb_tag_with_block_ram_1_io_raddr; // @[BTB.scala 249:54]
  wire [8:0] btb_tag_with_block_ram_1_io_waddr; // @[BTB.scala 249:54]
  wire [7:0] btb_tag_with_block_ram_1_io_wdata; // @[BTB.scala 249:54]
  wire [7:0] btb_tag_with_block_ram_1_io_rdata; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_2_clock; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_2_io_wen; // @[BTB.scala 249:54]
  wire [8:0] btb_tag_with_block_ram_2_io_raddr; // @[BTB.scala 249:54]
  wire [8:0] btb_tag_with_block_ram_2_io_waddr; // @[BTB.scala 249:54]
  wire [7:0] btb_tag_with_block_ram_2_io_wdata; // @[BTB.scala 249:54]
  wire [7:0] btb_tag_with_block_ram_2_io_rdata; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_3_clock; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_3_io_wen; // @[BTB.scala 249:54]
  wire [8:0] btb_tag_with_block_ram_3_io_raddr; // @[BTB.scala 249:54]
  wire [8:0] btb_tag_with_block_ram_3_io_waddr; // @[BTB.scala 249:54]
  wire [7:0] btb_tag_with_block_ram_3_io_wdata; // @[BTB.scala 249:54]
  wire [7:0] btb_tag_with_block_ram_3_io_rdata; // @[BTB.scala 249:54]
  wire  btb_data_with_block_ram_clock; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_io_wen; // @[BTB.scala 250:54]
  wire [8:0] btb_data_with_block_ram_io_raddr; // @[BTB.scala 250:54]
  wire [8:0] btb_data_with_block_ram_io_waddr; // @[BTB.scala 250:54]
  wire [31:0] btb_data_with_block_ram_io_wdata; // @[BTB.scala 250:54]
  wire [31:0] btb_data_with_block_ram_io_rdata; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_1_clock; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_1_io_wen; // @[BTB.scala 250:54]
  wire [8:0] btb_data_with_block_ram_1_io_raddr; // @[BTB.scala 250:54]
  wire [8:0] btb_data_with_block_ram_1_io_waddr; // @[BTB.scala 250:54]
  wire [31:0] btb_data_with_block_ram_1_io_wdata; // @[BTB.scala 250:54]
  wire [31:0] btb_data_with_block_ram_1_io_rdata; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_2_clock; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_2_io_wen; // @[BTB.scala 250:54]
  wire [8:0] btb_data_with_block_ram_2_io_raddr; // @[BTB.scala 250:54]
  wire [8:0] btb_data_with_block_ram_2_io_waddr; // @[BTB.scala 250:54]
  wire [31:0] btb_data_with_block_ram_2_io_wdata; // @[BTB.scala 250:54]
  wire [31:0] btb_data_with_block_ram_2_io_rdata; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_3_clock; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_3_io_wen; // @[BTB.scala 250:54]
  wire [8:0] btb_data_with_block_ram_3_io_raddr; // @[BTB.scala 250:54]
  wire [8:0] btb_data_with_block_ram_3_io_waddr; // @[BTB.scala 250:54]
  wire [31:0] btb_data_with_block_ram_3_io_wdata; // @[BTB.scala 250:54]
  wire [31:0] btb_data_with_block_ram_3_io_rdata; // @[BTB.scala 250:54]
  wire  _btb_banks_0_wen_T_1 = io_aw_addr[3:2] == 2'h0; // @[BTB.scala 253:62]
  wire  _btb_banks_1_wen_T_1 = io_aw_addr[3:2] == 2'h1; // @[BTB.scala 253:62]
  wire  _btb_banks_2_wen_T_1 = io_aw_addr[3:2] == 2'h2; // @[BTB.scala 253:62]
  wire  _btb_banks_3_wen_T_1 = io_aw_addr[3:2] == 2'h3; // @[BTB.scala 253:62]
  reg [31:0] ar_addr_reg; // @[BTB.scala 263:30]
  wire [31:0] btb_banks_0_rdata = btb_data_with_block_ram_io_rdata; // @[BTB.scala 250:{28,28}]
  wire [31:0] btb_banks_1_rdata = btb_data_with_block_ram_1_io_rdata; // @[BTB.scala 250:{28,28}]
  wire [31:0] _GEN_1 = 2'h1 == ar_addr_reg[3:2] ? btb_banks_1_rdata : btb_banks_0_rdata; // @[BTB.scala 265:{14,14}]
  wire [31:0] btb_banks_2_rdata = btb_data_with_block_ram_2_io_rdata; // @[BTB.scala 250:{28,28}]
  wire [31:0] _GEN_2 = 2'h2 == ar_addr_reg[3:2] ? btb_banks_2_rdata : _GEN_1; // @[BTB.scala 265:{14,14}]
  wire [31:0] btb_banks_3_rdata = btb_data_with_block_ram_3_io_rdata; // @[BTB.scala 250:{28,28}]
  wire [4:0] _tag_banks_0_wdata_T_1 = {1'h1,io_aw_addr[16:13]}; // @[Cat.scala 31:58]
  wire [7:0] tag_banks_0_rdata = btb_tag_with_block_ram_io_rdata; // @[BTB.scala 249:{28,28}]
  wire [7:0] tag_banks_1_rdata = btb_tag_with_block_ram_1_io_rdata; // @[BTB.scala 249:{28,28}]
  wire [7:0] _GEN_13 = 2'h1 == ar_addr_reg[3:2] ? tag_banks_1_rdata : tag_banks_0_rdata; // @[BTB.scala 286:{67,67}]
  wire [7:0] tag_banks_2_rdata = btb_tag_with_block_ram_2_io_rdata; // @[BTB.scala 249:{28,28}]
  wire [7:0] _GEN_14 = 2'h2 == ar_addr_reg[3:2] ? tag_banks_2_rdata : _GEN_13; // @[BTB.scala 286:{67,67}]
  wire [7:0] tag_banks_3_rdata = btb_tag_with_block_ram_3_io_rdata; // @[BTB.scala 249:{28,28}]
  wire [7:0] _GEN_15 = 2'h3 == ar_addr_reg[3:2] ? tag_banks_3_rdata : _GEN_14; // @[BTB.scala 286:{67,67}]
  btb_tag_with_block_ram btb_tag_with_block_ram ( // @[BTB.scala 249:54]
    .clock(btb_tag_with_block_ram_clock),
    .io_wen(btb_tag_with_block_ram_io_wen),
    .io_raddr(btb_tag_with_block_ram_io_raddr),
    .io_waddr(btb_tag_with_block_ram_io_waddr),
    .io_wdata(btb_tag_with_block_ram_io_wdata),
    .io_rdata(btb_tag_with_block_ram_io_rdata)
  );
  btb_tag_with_block_ram btb_tag_with_block_ram_1 ( // @[BTB.scala 249:54]
    .clock(btb_tag_with_block_ram_1_clock),
    .io_wen(btb_tag_with_block_ram_1_io_wen),
    .io_raddr(btb_tag_with_block_ram_1_io_raddr),
    .io_waddr(btb_tag_with_block_ram_1_io_waddr),
    .io_wdata(btb_tag_with_block_ram_1_io_wdata),
    .io_rdata(btb_tag_with_block_ram_1_io_rdata)
  );
  btb_tag_with_block_ram btb_tag_with_block_ram_2 ( // @[BTB.scala 249:54]
    .clock(btb_tag_with_block_ram_2_clock),
    .io_wen(btb_tag_with_block_ram_2_io_wen),
    .io_raddr(btb_tag_with_block_ram_2_io_raddr),
    .io_waddr(btb_tag_with_block_ram_2_io_waddr),
    .io_wdata(btb_tag_with_block_ram_2_io_wdata),
    .io_rdata(btb_tag_with_block_ram_2_io_rdata)
  );
  btb_tag_with_block_ram btb_tag_with_block_ram_3 ( // @[BTB.scala 249:54]
    .clock(btb_tag_with_block_ram_3_clock),
    .io_wen(btb_tag_with_block_ram_3_io_wen),
    .io_raddr(btb_tag_with_block_ram_3_io_raddr),
    .io_waddr(btb_tag_with_block_ram_3_io_waddr),
    .io_wdata(btb_tag_with_block_ram_3_io_wdata),
    .io_rdata(btb_tag_with_block_ram_3_io_rdata)
  );
  btb_data_with_block_ram btb_data_with_block_ram ( // @[BTB.scala 250:54]
    .clock(btb_data_with_block_ram_clock),
    .io_wen(btb_data_with_block_ram_io_wen),
    .io_raddr(btb_data_with_block_ram_io_raddr),
    .io_waddr(btb_data_with_block_ram_io_waddr),
    .io_wdata(btb_data_with_block_ram_io_wdata),
    .io_rdata(btb_data_with_block_ram_io_rdata)
  );
  btb_data_with_block_ram btb_data_with_block_ram_1 ( // @[BTB.scala 250:54]
    .clock(btb_data_with_block_ram_1_clock),
    .io_wen(btb_data_with_block_ram_1_io_wen),
    .io_raddr(btb_data_with_block_ram_1_io_raddr),
    .io_waddr(btb_data_with_block_ram_1_io_waddr),
    .io_wdata(btb_data_with_block_ram_1_io_wdata),
    .io_rdata(btb_data_with_block_ram_1_io_rdata)
  );
  btb_data_with_block_ram btb_data_with_block_ram_2 ( // @[BTB.scala 250:54]
    .clock(btb_data_with_block_ram_2_clock),
    .io_wen(btb_data_with_block_ram_2_io_wen),
    .io_raddr(btb_data_with_block_ram_2_io_raddr),
    .io_waddr(btb_data_with_block_ram_2_io_waddr),
    .io_wdata(btb_data_with_block_ram_2_io_wdata),
    .io_rdata(btb_data_with_block_ram_2_io_rdata)
  );
  btb_data_with_block_ram btb_data_with_block_ram_3 ( // @[BTB.scala 250:54]
    .clock(btb_data_with_block_ram_3_clock),
    .io_wen(btb_data_with_block_ram_3_io_wen),
    .io_raddr(btb_data_with_block_ram_3_io_raddr),
    .io_waddr(btb_data_with_block_ram_3_io_waddr),
    .io_wdata(btb_data_with_block_ram_3_io_wdata),
    .io_rdata(btb_data_with_block_ram_3_io_rdata)
  );
  assign io_out_L = 2'h3 == ar_addr_reg[3:2] ? btb_banks_3_rdata : _GEN_2; // @[BTB.scala 265:{14,14}]
  assign io_hit_L = _GEN_15[3:0] == io_ar_addr_L[16:13] & _GEN_15[4]; // @[BTB.scala 286:167]
  assign btb_tag_with_block_ram_clock = clock;
  assign btb_tag_with_block_ram_io_wen = _btb_banks_0_wen_T_1 & io_write; // @[BTB.scala 271:75]
  assign btb_tag_with_block_ram_io_raddr = io_ar_addr_L[12:4]; // @[BTB.scala 273:43]
  assign btb_tag_with_block_ram_io_waddr = io_aw_addr[12:4]; // @[BTB.scala 279:41]
  assign btb_tag_with_block_ram_io_wdata = {{3'd0}, _tag_banks_0_wdata_T_1}; // @[BTB.scala 249:28 272:28]
  assign btb_tag_with_block_ram_1_clock = clock;
  assign btb_tag_with_block_ram_1_io_wen = _btb_banks_1_wen_T_1 & io_write; // @[BTB.scala 271:75]
  assign btb_tag_with_block_ram_1_io_raddr = io_ar_addr_L[12:4]; // @[BTB.scala 273:43]
  assign btb_tag_with_block_ram_1_io_waddr = io_aw_addr[12:4]; // @[BTB.scala 279:41]
  assign btb_tag_with_block_ram_1_io_wdata = {{3'd0}, _tag_banks_0_wdata_T_1}; // @[BTB.scala 249:28 272:28]
  assign btb_tag_with_block_ram_2_clock = clock;
  assign btb_tag_with_block_ram_2_io_wen = _btb_banks_2_wen_T_1 & io_write; // @[BTB.scala 271:75]
  assign btb_tag_with_block_ram_2_io_raddr = io_ar_addr_L[12:4]; // @[BTB.scala 273:43]
  assign btb_tag_with_block_ram_2_io_waddr = io_aw_addr[12:4]; // @[BTB.scala 279:41]
  assign btb_tag_with_block_ram_2_io_wdata = {{3'd0}, _tag_banks_0_wdata_T_1}; // @[BTB.scala 249:28 272:28]
  assign btb_tag_with_block_ram_3_clock = clock;
  assign btb_tag_with_block_ram_3_io_wen = _btb_banks_3_wen_T_1 & io_write; // @[BTB.scala 271:75]
  assign btb_tag_with_block_ram_3_io_raddr = io_ar_addr_L[12:4]; // @[BTB.scala 273:43]
  assign btb_tag_with_block_ram_3_io_waddr = io_aw_addr[12:4]; // @[BTB.scala 279:41]
  assign btb_tag_with_block_ram_3_io_wdata = {{3'd0}, _tag_banks_0_wdata_T_1}; // @[BTB.scala 249:28 272:28]
  assign btb_data_with_block_ram_clock = clock;
  assign btb_data_with_block_ram_io_wen = io_aw_addr[3:2] == 2'h0 & io_write; // @[BTB.scala 253:75]
  assign btb_data_with_block_ram_io_raddr = io_ar_addr_L[12:4]; // @[BTB.scala 255:43]
  assign btb_data_with_block_ram_io_waddr = io_aw_addr[12:4]; // @[BTB.scala 261:41]
  assign btb_data_with_block_ram_io_wdata = io_aw_target_addr; // @[BTB.scala 250:28 254:28]
  assign btb_data_with_block_ram_1_clock = clock;
  assign btb_data_with_block_ram_1_io_wen = io_aw_addr[3:2] == 2'h1 & io_write; // @[BTB.scala 253:75]
  assign btb_data_with_block_ram_1_io_raddr = io_ar_addr_L[12:4]; // @[BTB.scala 255:43]
  assign btb_data_with_block_ram_1_io_waddr = io_aw_addr[12:4]; // @[BTB.scala 261:41]
  assign btb_data_with_block_ram_1_io_wdata = io_aw_target_addr; // @[BTB.scala 250:28 254:28]
  assign btb_data_with_block_ram_2_clock = clock;
  assign btb_data_with_block_ram_2_io_wen = io_aw_addr[3:2] == 2'h2 & io_write; // @[BTB.scala 253:75]
  assign btb_data_with_block_ram_2_io_raddr = io_ar_addr_L[12:4]; // @[BTB.scala 255:43]
  assign btb_data_with_block_ram_2_io_waddr = io_aw_addr[12:4]; // @[BTB.scala 261:41]
  assign btb_data_with_block_ram_2_io_wdata = io_aw_target_addr; // @[BTB.scala 250:28 254:28]
  assign btb_data_with_block_ram_3_clock = clock;
  assign btb_data_with_block_ram_3_io_wen = io_aw_addr[3:2] == 2'h3 & io_write; // @[BTB.scala 253:75]
  assign btb_data_with_block_ram_3_io_raddr = io_ar_addr_L[12:4]; // @[BTB.scala 255:43]
  assign btb_data_with_block_ram_3_io_waddr = io_aw_addr[12:4]; // @[BTB.scala 261:41]
  assign btb_data_with_block_ram_3_io_wdata = io_aw_target_addr; // @[BTB.scala 250:28 254:28]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BTB.scala 263:30]
      ar_addr_reg <= 32'h0; // @[BTB.scala 263:30]
    end else begin
      ar_addr_reg <= io_ar_addr_L; // @[BTB.scala 264:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ar_addr_reg = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    ar_addr_reg = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module branch_prediction_with_blockram(
  input         clock,
  input         reset,
  input  [31:0] io_pc,
  input  [31:0] io_write_pc,
  input  [3:0]  io_aw_pht_ways_addr,
  input  [6:0]  io_aw_pht_addr,
  input  [6:0]  io_aw_bht_addr,
  input  [31:0] io_aw_target_addr,
  input         io_btb_write,
  input         io_bht_write,
  input         io_pht_write,
  input  [6:0]  io_bht_in,
  input  [7:0]  io_pht_in,
  output [1:0]  io_out_L,
  output        io_pre_L,
  output [6:0]  io_bht_L,
  output        io_btb_hit_0,
  output [31:0] io_pre_target_L,
  input         io_stage2_stall,
  input         io_stage2_flush,
  output [7:0]  io_pht_out,
  output [6:0]  io_lookup_data_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  PHTS_banks_oneissue_block_ram_clock; // @[branch_prediction.scala 200:28]
  wire  PHTS_banks_oneissue_block_ram_reset; // @[branch_prediction.scala 200:28]
  wire [1:0] PHTS_banks_oneissue_block_ram_io_ar_bank_sel; // @[branch_prediction.scala 200:28]
  wire [6:0] PHTS_banks_oneissue_block_ram_io_ar_addr_L; // @[branch_prediction.scala 200:28]
  wire [2:0] PHTS_banks_oneissue_block_ram_io_ar_pht_addr; // @[branch_prediction.scala 200:28]
  wire [6:0] PHTS_banks_oneissue_block_ram_io_aw_addr; // @[branch_prediction.scala 200:28]
  wire [2:0] PHTS_banks_oneissue_block_ram_io_aw_pht_addr; // @[branch_prediction.scala 200:28]
  wire [1:0] PHTS_banks_oneissue_block_ram_io_aw_bank_sel; // @[branch_prediction.scala 200:28]
  wire  PHTS_banks_oneissue_block_ram_io_write; // @[branch_prediction.scala 200:28]
  wire [7:0] PHTS_banks_oneissue_block_ram_io_in; // @[branch_prediction.scala 200:28]
  wire [1:0] PHTS_banks_oneissue_block_ram_io_out_L; // @[branch_prediction.scala 200:28]
  wire [7:0] PHTS_banks_oneissue_block_ram_io_pht_out; // @[branch_prediction.scala 200:28]
  wire  BHT_banks_oneissue_clock; // @[branch_prediction.scala 201:28]
  wire  BHT_banks_oneissue_reset; // @[branch_prediction.scala 201:28]
  wire [1:0] BHT_banks_oneissue_io_ar_bank_sel; // @[branch_prediction.scala 201:28]
  wire [6:0] BHT_banks_oneissue_io_ar_addr_L; // @[branch_prediction.scala 201:28]
  wire [6:0] BHT_banks_oneissue_io_aw_addr; // @[branch_prediction.scala 201:28]
  wire  BHT_banks_oneissue_io_write; // @[branch_prediction.scala 201:28]
  wire [2:0] BHT_banks_oneissue_io_in; // @[branch_prediction.scala 201:28]
  wire [2:0] BHT_banks_oneissue_io_out_L; // @[branch_prediction.scala 201:28]
  wire  BTB_banks_oneissue_with_block_ram_clock; // @[branch_prediction.scala 202:27]
  wire  BTB_banks_oneissue_with_block_ram_reset; // @[branch_prediction.scala 202:27]
  wire [31:0] BTB_banks_oneissue_with_block_ram_io_ar_addr_L; // @[branch_prediction.scala 202:27]
  wire [31:0] BTB_banks_oneissue_with_block_ram_io_aw_addr; // @[branch_prediction.scala 202:27]
  wire [31:0] BTB_banks_oneissue_with_block_ram_io_aw_target_addr; // @[branch_prediction.scala 202:27]
  wire  BTB_banks_oneissue_with_block_ram_io_write; // @[branch_prediction.scala 202:27]
  wire [31:0] BTB_banks_oneissue_with_block_ram_io_out_L; // @[branch_prediction.scala 202:27]
  wire  BTB_banks_oneissue_with_block_ram_io_hit_L; // @[branch_prediction.scala 202:27]
  wire  pc_hash_num_array_0 = ^io_pc[7:4]; // @[macros.scala 389:45]
  wire  pc_hash_num_array_1 = ^io_pc[11:8]; // @[macros.scala 389:45]
  wire  pc_hash_num_array_2 = ^io_pc[15:12]; // @[macros.scala 389:45]
  wire  pc_hash_num_array_3 = ^io_pc[19:16]; // @[macros.scala 389:45]
  wire [3:0] pc_hash = {pc_hash_num_array_3,pc_hash_num_array_2,pc_hash_num_array_1,pc_hash_num_array_0}; // @[macros.scala 391:13]
  reg [6:0] stage_2_pht_lookup_0; // @[branch_prediction.scala 204:37]
  wire [6:0] stage_1_pht_lookup_0 = {BHT_banks_oneissue_io_out_L,io_pc[14:11]}; // @[Cat.scala 31:58]
  wire  _io_pre_L_T_1 = 2'h0 == io_out_L ? 1'h0 : 1'h1; // @[Mux.scala 81:58]
  wire  _io_pre_L_T_3 = 2'h1 == io_out_L ? 1'h0 : _io_pre_L_T_1; // @[Mux.scala 81:58]
  PHTS_banks_oneissue_block_ram PHTS_banks_oneissue_block_ram ( // @[branch_prediction.scala 200:28]
    .clock(PHTS_banks_oneissue_block_ram_clock),
    .reset(PHTS_banks_oneissue_block_ram_reset),
    .io_ar_bank_sel(PHTS_banks_oneissue_block_ram_io_ar_bank_sel),
    .io_ar_addr_L(PHTS_banks_oneissue_block_ram_io_ar_addr_L),
    .io_ar_pht_addr(PHTS_banks_oneissue_block_ram_io_ar_pht_addr),
    .io_aw_addr(PHTS_banks_oneissue_block_ram_io_aw_addr),
    .io_aw_pht_addr(PHTS_banks_oneissue_block_ram_io_aw_pht_addr),
    .io_aw_bank_sel(PHTS_banks_oneissue_block_ram_io_aw_bank_sel),
    .io_write(PHTS_banks_oneissue_block_ram_io_write),
    .io_in(PHTS_banks_oneissue_block_ram_io_in),
    .io_out_L(PHTS_banks_oneissue_block_ram_io_out_L),
    .io_pht_out(PHTS_banks_oneissue_block_ram_io_pht_out)
  );
  BHT_banks_oneissue BHT_banks_oneissue ( // @[branch_prediction.scala 201:28]
    .clock(BHT_banks_oneissue_clock),
    .reset(BHT_banks_oneissue_reset),
    .io_ar_bank_sel(BHT_banks_oneissue_io_ar_bank_sel),
    .io_ar_addr_L(BHT_banks_oneissue_io_ar_addr_L),
    .io_aw_addr(BHT_banks_oneissue_io_aw_addr),
    .io_write(BHT_banks_oneissue_io_write),
    .io_in(BHT_banks_oneissue_io_in),
    .io_out_L(BHT_banks_oneissue_io_out_L)
  );
  BTB_banks_oneissue_with_block_ram BTB_banks_oneissue_with_block_ram ( // @[branch_prediction.scala 202:27]
    .clock(BTB_banks_oneissue_with_block_ram_clock),
    .reset(BTB_banks_oneissue_with_block_ram_reset),
    .io_ar_addr_L(BTB_banks_oneissue_with_block_ram_io_ar_addr_L),
    .io_aw_addr(BTB_banks_oneissue_with_block_ram_io_aw_addr),
    .io_aw_target_addr(BTB_banks_oneissue_with_block_ram_io_aw_target_addr),
    .io_write(BTB_banks_oneissue_with_block_ram_io_write),
    .io_out_L(BTB_banks_oneissue_with_block_ram_io_out_L),
    .io_hit_L(BTB_banks_oneissue_with_block_ram_io_hit_L)
  );
  assign io_out_L = PHTS_banks_oneissue_block_ram_io_out_L; // @[branch_prediction.scala 286:14]
  assign io_pre_L = 2'h2 == io_out_L | _io_pre_L_T_3; // @[Mux.scala 81:58]
  assign io_bht_L = {{4'd0}, BHT_banks_oneissue_io_out_L}; // @[branch_prediction.scala 290:14]
  assign io_btb_hit_0 = BTB_banks_oneissue_with_block_ram_io_hit_L; // @[branch_prediction.scala 302:19]
  assign io_pre_target_L = BTB_banks_oneissue_with_block_ram_io_out_L; // @[branch_prediction.scala 298:21]
  assign io_pht_out = PHTS_banks_oneissue_block_ram_io_pht_out; // @[branch_prediction.scala 306:16]
  assign io_lookup_data_0 = stage_2_pht_lookup_0; // @[branch_prediction.scala 229:23]
  assign PHTS_banks_oneissue_block_ram_clock = clock;
  assign PHTS_banks_oneissue_block_ram_reset = reset;
  assign PHTS_banks_oneissue_block_ram_io_ar_bank_sel = io_pc[3:2]; // @[branch_prediction.scala 243:36]
  assign PHTS_banks_oneissue_block_ram_io_ar_addr_L = {BHT_banks_oneissue_io_out_L,io_pc[14:11]}; // @[Cat.scala 31:58]
  assign PHTS_banks_oneissue_block_ram_io_ar_pht_addr = pc_hash[2:0]; // @[branch_prediction.scala 244:28]
  assign PHTS_banks_oneissue_block_ram_io_aw_addr = io_aw_pht_addr; // @[branch_prediction.scala 259:24]
  assign PHTS_banks_oneissue_block_ram_io_aw_pht_addr = io_aw_pht_ways_addr[2:0]; // @[branch_prediction.scala 260:28]
  assign PHTS_banks_oneissue_block_ram_io_aw_bank_sel = io_write_pc[3:2]; // @[branch_prediction.scala 261:42]
  assign PHTS_banks_oneissue_block_ram_io_write = io_pht_write; // @[branch_prediction.scala 262:22]
  assign PHTS_banks_oneissue_block_ram_io_in = io_pht_in; // @[branch_prediction.scala 263:19]
  assign BHT_banks_oneissue_clock = clock;
  assign BHT_banks_oneissue_reset = reset;
  assign BHT_banks_oneissue_io_ar_bank_sel = io_pc[3:2]; // @[branch_prediction.scala 235:36]
  assign BHT_banks_oneissue_io_ar_addr_L = io_pc[10:4]; // @[branch_prediction.scala 237:34]
  assign BHT_banks_oneissue_io_aw_addr = io_aw_bht_addr; // @[branch_prediction.scala 241:24]
  assign BHT_banks_oneissue_io_write = io_bht_write; // @[branch_prediction.scala 236:22]
  assign BHT_banks_oneissue_io_in = io_bht_in[2:0]; // @[branch_prediction.scala 240:19]
  assign BTB_banks_oneissue_with_block_ram_clock = clock;
  assign BTB_banks_oneissue_with_block_ram_reset = reset;
  assign BTB_banks_oneissue_with_block_ram_io_ar_addr_L = io_pc; // @[branch_prediction.scala 266:25]
  assign BTB_banks_oneissue_with_block_ram_io_aw_addr = io_write_pc; // @[branch_prediction.scala 269:25]
  assign BTB_banks_oneissue_with_block_ram_io_aw_target_addr = io_aw_target_addr; // @[branch_prediction.scala 270:30]
  assign BTB_banks_oneissue_with_block_ram_io_write = io_btb_write; // @[branch_prediction.scala 271:21]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[branch_prediction.scala 218:33]
      stage_2_pht_lookup_0 <= 7'h0;
    end else if (io_stage2_flush) begin // @[branch_prediction.scala 218:57]
      stage_2_pht_lookup_0 <= 7'h0;
    end else if (io_stage2_stall) begin
      stage_2_pht_lookup_0 <= stage_1_pht_lookup_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stage_2_pht_lookup_0 = _RAND_0[6:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    stage_2_pht_lookup_0 = 7'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module bru_detail(
  input         clock,
  input         reset,
  input         io_stall,
  input         io_flush,
  input  [1:0]  io_in_pht,
  input  [6:0]  io_in_bht,
  input  [3:0]  io_in_hashcode,
  input  [31:0] io_in_target_pc,
  input  [6:0]  io_in_lookup_data,
  input  [7:0]  io_in_pht_lookup_value,
  output [1:0]  io_out_pht,
  output [6:0]  io_out_bht,
  output [3:0]  io_out_hashcode,
  output [31:0] io_out_target_pc,
  output [6:0]  io_out_lookup_data,
  output [7:0]  io_out_pht_lookup_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] pht_value; // @[myCPU.scala 625:30]
  reg [6:0] bht_value; // @[myCPU.scala 626:30]
  reg [3:0] hashcode_value; // @[myCPU.scala 627:35]
  reg [31:0] target_pc_value; // @[myCPU.scala 628:36]
  reg [6:0] lookup_data_value; // @[myCPU.scala 629:38]
  reg [7:0] pht_lookup_value_data; // @[myCPU.scala 630:42]
  assign io_out_pht = pht_value; // @[myCPU.scala 639:16]
  assign io_out_bht = bht_value; // @[myCPU.scala 640:16]
  assign io_out_hashcode = hashcode_value; // @[myCPU.scala 641:21]
  assign io_out_target_pc = target_pc_value; // @[myCPU.scala 642:22]
  assign io_out_lookup_data = lookup_data_value; // @[myCPU.scala 643:24]
  assign io_out_pht_lookup_value = pht_lookup_value_data; // @[myCPU.scala 644:29]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[myCPU.scala 631:21]
      pht_value <= 2'h0;
    end else if (io_flush) begin // @[myCPU.scala 631:38]
      pht_value <= 2'h0;
    end else if (io_stall) begin
      pht_value <= io_in_pht;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[myCPU.scala 632:21]
      bht_value <= 7'h0;
    end else if (io_flush) begin // @[myCPU.scala 632:38]
      bht_value <= 7'h0;
    end else if (io_stall) begin
      bht_value <= io_in_bht;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[myCPU.scala 633:26]
      hashcode_value <= 4'h0;
    end else if (io_flush) begin // @[myCPU.scala 633:43]
      hashcode_value <= 4'h0;
    end else if (io_stall) begin
      hashcode_value <= io_in_hashcode;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[myCPU.scala 634:27]
      target_pc_value <= 32'h0;
    end else if (io_flush) begin // @[myCPU.scala 634:44]
      target_pc_value <= 32'h0;
    end else if (io_stall) begin
      target_pc_value <= io_in_target_pc;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[myCPU.scala 635:29]
      lookup_data_value <= 7'h0;
    end else if (io_flush) begin // @[myCPU.scala 635:46]
      lookup_data_value <= 7'h0;
    end else if (io_stall) begin
      lookup_data_value <= io_in_lookup_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[myCPU.scala 636:33]
      pht_lookup_value_data <= 8'h0;
    end else if (io_flush) begin // @[myCPU.scala 636:50]
      pht_lookup_value_data <= 8'h0;
    end else if (io_stall) begin
      pht_lookup_value_data <= io_in_pht_lookup_value;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pht_value = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  bht_value = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  hashcode_value = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  target_pc_value = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  lookup_data_value = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  pht_lookup_value_data = _RAND_5[7:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    pht_value = 2'h0;
  end
  if (reset) begin
    bht_value = 7'h0;
  end
  if (reset) begin
    hashcode_value = 4'h0;
  end
  if (reset) begin
    target_pc_value = 32'h0;
  end
  if (reset) begin
    lookup_data_value = 7'h0;
  end
  if (reset) begin
    pht_lookup_value_data = 8'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module tlb_data_register(
  input         clock,
  input         reset,
  input         io_flush,
  input         io_stall,
  output [18:0] io_tlb_read_data_vaddr,
  output [7:0]  io_tlb_read_data_asid,
  output        io_tlb_read_data_g,
  output [19:0] io_tlb_read_data_paddr_0,
  output [19:0] io_tlb_read_data_paddr_1,
  output [2:0]  io_tlb_read_data_c_0,
  output [2:0]  io_tlb_read_data_c_1,
  output        io_tlb_read_data_d_0,
  output        io_tlb_read_data_d_1,
  output        io_tlb_read_data_v_0,
  output        io_tlb_read_data_v_1,
  input  [18:0] io_tlb_write_data_vaddr,
  input  [7:0]  io_tlb_write_data_asid,
  input         io_tlb_write_data_g,
  input  [19:0] io_tlb_write_data_paddr_0,
  input  [19:0] io_tlb_write_data_paddr_1,
  input  [2:0]  io_tlb_write_data_c_0,
  input  [2:0]  io_tlb_write_data_c_1,
  input         io_tlb_write_data_d_0,
  input         io_tlb_write_data_d_1,
  input         io_tlb_write_data_v_0,
  input         io_tlb_write_data_v_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [77:0] tlb_data_reg; // @[myCPU.scala 952:31]
  wire [25:0] tlb_data_reg_lo = {io_tlb_write_data_v_0,io_tlb_write_data_paddr_1,io_tlb_write_data_c_1,
    io_tlb_write_data_d_1,io_tlb_write_data_v_1}; // @[Cat.scala 31:58]
  wire [77:0] _tlb_data_reg_T = {io_tlb_write_data_vaddr,io_tlb_write_data_asid,io_tlb_write_data_g,
    io_tlb_write_data_paddr_0,io_tlb_write_data_c_0,io_tlb_write_data_d_0,tlb_data_reg_lo}; // @[Cat.scala 31:58]
  assign io_tlb_read_data_vaddr = tlb_data_reg[77:59]; // @[macros.scala 432:43]
  assign io_tlb_read_data_asid = tlb_data_reg[58:51]; // @[macros.scala 431:43]
  assign io_tlb_read_data_g = tlb_data_reg[50]; // @[macros.scala 430:41]
  assign io_tlb_read_data_paddr_0 = tlb_data_reg[49:30]; // @[macros.scala 429:47]
  assign io_tlb_read_data_paddr_1 = tlb_data_reg[24:5]; // @[macros.scala 427:47]
  assign io_tlb_read_data_c_0 = tlb_data_reg[29:27]; // @[myCPU.scala 959:56]
  assign io_tlb_read_data_c_1 = tlb_data_reg[4:2]; // @[myCPU.scala 956:56]
  assign io_tlb_read_data_d_0 = tlb_data_reg[26]; // @[myCPU.scala 958:56]
  assign io_tlb_read_data_d_1 = tlb_data_reg[1]; // @[myCPU.scala 955:56]
  assign io_tlb_read_data_v_0 = tlb_data_reg[25]; // @[myCPU.scala 957:56]
  assign io_tlb_read_data_v_1 = tlb_data_reg[0]; // @[myCPU.scala 954:56]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[myCPU.scala 953:24]
      tlb_data_reg <= 78'h0;
    end else if (io_flush) begin // @[myCPU.scala 953:41]
      tlb_data_reg <= 78'h0;
    end else if (io_stall) begin
      tlb_data_reg <= _tlb_data_reg_T;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  tlb_data_reg = _RAND_0[77:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    tlb_data_reg = 78'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module myCPU(
  input  [5:0]  ext_int,
  input         resetn,
  input         clk,
  output        inst_cache,
  output        inst_sram_en,
  output [31:0] inst_sram_addr,
  input  [39:0] inst_sram_rdata_L,
  input  [1:0]  inst_write_en,
  output        inst_ready_branch,
  output        inst_buffer_empty,
  output [7:0]  cp0_asid,
  input  [1:0]  inst_tlb_exception,
  output        stage2_flush,
  input         stage2_stall,
  output [1:0]  stage1_valid_flush,
  output        inst_ready_to_use,
  output        inst_buffer_full,
  output        data_sram_en,
  output        data_sram_wen,
  output [1:0]  data_size,
  output [31:0] data_sram_addr,
  output [31:0] data_sram_wdata,
  output        data_cache,
  input  [31:0] data_sram_rdata,
  input         data_stage2_stall,
  input  [2:0]  data_tlb_exception,
  output [3:0]  data_wstrb,
  output [31:0] tlbp_search_vaddr,
  output        tlbp_search_en,
  input  [3:0]  tlb_search_index,
  input         tlb_search_hit,
  output [3:0]  tlb_read_index,
  output [3:0]  tlb_write_index,
  output [31:0] debug_wb_pc,
  output [3:0]  debug_wb_rf_wen,
  output [4:0]  debug_wb_rf_wnum,
  output [31:0] debug_wb_rf_wdata,
  output [18:0] cp0_tlb_read_data_vaddr,
  output [7:0]  cp0_tlb_read_data_asid,
  output        cp0_tlb_read_data_g,
  output [19:0] cp0_tlb_read_data_paddr_0,
  output [19:0] cp0_tlb_read_data_paddr_1,
  output [2:0]  cp0_tlb_read_data_c_0,
  output [2:0]  cp0_tlb_read_data_c_1,
  output        cp0_tlb_read_data_d_0,
  output        cp0_tlb_read_data_d_1,
  output        cp0_tlb_read_data_v_0,
  output        cp0_tlb_read_data_v_1,
  input  [18:0] cp0_tlb_write_data_vaddr,
  input  [7:0]  cp0_tlb_write_data_asid,
  input         cp0_tlb_write_data_g,
  input  [19:0] cp0_tlb_write_data_paddr_0,
  input  [19:0] cp0_tlb_write_data_paddr_1,
  input  [2:0]  cp0_tlb_write_data_c_0,
  input  [2:0]  cp0_tlb_write_data_c_1,
  input         cp0_tlb_write_data_d_0,
  input         cp0_tlb_write_data_d_1,
  input         cp0_tlb_write_data_v_0,
  input         cp0_tlb_write_data_v_1,
  output        tlb_write_en
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
`endif // RANDOMIZE_REG_INIT
  wire [23:0] _alu_io_ctrl; // @[myCPU.scala 120:22]
  wire [31:0] _alu_io_in1; // @[myCPU.scala 120:22]
  wire [31:0] _alu_io_in2; // @[myCPU.scala 120:22]
  wire [31:0] _alu_io_result; // @[myCPU.scala 120:22]
  wire  _alu_io_overflow; // @[myCPU.scala 120:22]
  wire  _br_reset; // @[myCPU.scala 121:22]
  wire [31:0] _br_io_rs; // @[myCPU.scala 121:22]
  wire [31:0] _br_io_rt; // @[myCPU.scala 121:22]
  wire [5:0] _br_io_branch; // @[myCPU.scala 121:22]
  wire  _br_io_exe; // @[myCPU.scala 121:22]
  wire  _cfu_reset; // @[myCPU.scala 122:22]
  wire  _cfu_io_Inst_Fifo_Empty; // @[myCPU.scala 122:22]
  wire  _cfu_io_dmem_calD; // @[myCPU.scala 122:22]
  wire  _cfu_io_BranchD_Flag; // @[myCPU.scala 122:22]
  wire  _cfu_io_JRD; // @[myCPU.scala 122:22]
  wire  _cfu_io_CanBranchD; // @[myCPU.scala 122:22]
  wire  _cfu_io_DivPendingE; // @[myCPU.scala 122:22]
  wire  _cfu_io_DataPendingM; // @[myCPU.scala 122:22]
  wire  _cfu_io_InException; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_WriteRegE; // @[myCPU.scala 122:22]
  wire  _cfu_io_RegWriteE; // @[myCPU.scala 122:22]
  wire [1:0] _cfu_io_HiLoToRegE; // @[myCPU.scala 122:22]
  wire  _cfu_io_CP0ToRegE; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_WriteRegM; // @[myCPU.scala 122:22]
  wire  _cfu_io_MemToRegM; // @[myCPU.scala 122:22]
  wire  _cfu_io_RegWriteM; // @[myCPU.scala 122:22]
  wire [1:0] _cfu_io_HiLoWriteM; // @[myCPU.scala 122:22]
  wire  _cfu_io_CP0WriteM; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_WriteRegM2; // @[myCPU.scala 122:22]
  wire  _cfu_io_MemToRegM2; // @[myCPU.scala 122:22]
  wire  _cfu_io_RegWriteM2; // @[myCPU.scala 122:22]
  wire [1:0] _cfu_io_HiLoWriteM2; // @[myCPU.scala 122:22]
  wire  _cfu_io_CP0WriteM2; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_WriteRegW; // @[myCPU.scala 122:22]
  wire  _cfu_io_RegWriteW; // @[myCPU.scala 122:22]
  wire [1:0] _cfu_io_HiLoWriteW; // @[myCPU.scala 122:22]
  wire  _cfu_io_CP0WriteW; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_ReadCP0AddrE; // @[myCPU.scala 122:22]
  wire [2:0] _cfu_io_ReadCP0SelE; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_WriteCP0AddrM; // @[myCPU.scala 122:22]
  wire [2:0] _cfu_io_WriteCP0SelM; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_WriteCP0AddrM2; // @[myCPU.scala 122:22]
  wire [2:0] _cfu_io_WriteCP0SelM2; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_RsD; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_RtD; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_RsE; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_RtE; // @[myCPU.scala 122:22]
  wire  _cfu_io_StallF; // @[myCPU.scala 122:22]
  wire  _cfu_io_StallD; // @[myCPU.scala 122:22]
  wire  _cfu_io_StallE; // @[myCPU.scala 122:22]
  wire  _cfu_io_StallM; // @[myCPU.scala 122:22]
  wire  _cfu_io_StallM2; // @[myCPU.scala 122:22]
  wire  _cfu_io_StallW; // @[myCPU.scala 122:22]
  wire  _cfu_io_FlushD; // @[myCPU.scala 122:22]
  wire  _cfu_io_FlushE; // @[myCPU.scala 122:22]
  wire  _cfu_io_FlushM; // @[myCPU.scala 122:22]
  wire  _cfu_io_FlushM2; // @[myCPU.scala 122:22]
  wire  _cfu_io_FlushW; // @[myCPU.scala 122:22]
  wire [1:0] _cfu_io_ForwardAE; // @[myCPU.scala 122:22]
  wire [1:0] _cfu_io_ForwardBE; // @[myCPU.scala 122:22]
  wire [1:0] _cfu_io_ForwardAD; // @[myCPU.scala 122:22]
  wire [1:0] _cfu_io_ForwardBD; // @[myCPU.scala 122:22]
  wire [1:0] _cfu_io_ForwardHE; // @[myCPU.scala 122:22]
  wire [1:0] _cfu_io_ForwardCP0E; // @[myCPU.scala 122:22]
  wire  _cp0_clock; // @[myCPU.scala 123:22]
  wire  _cp0_reset; // @[myCPU.scala 123:22]
  wire [4:0] _cp0_io_cp0_read_addr; // @[myCPU.scala 123:22]
  wire [2:0] _cp0_io_cp0_read_sel; // @[myCPU.scala 123:22]
  wire [4:0] _cp0_io_cp0_write_addr; // @[myCPU.scala 123:22]
  wire [2:0] _cp0_io_cp0_write_sel; // @[myCPU.scala 123:22]
  wire [31:0] _cp0_io_cp0_write_data; // @[myCPU.scala 123:22]
  wire  _cp0_io_cp0_write_en; // @[myCPU.scala 123:22]
  wire [5:0] _cp0_io_int_i; // @[myCPU.scala 123:22]
  wire  _cp0_io_timer_int_has; // @[myCPU.scala 123:22]
  wire [31:0] _cp0_io_pc; // @[myCPU.scala 123:22]
  wire [31:0] _cp0_io_mem_bad_vaddr; // @[myCPU.scala 123:22]
  wire [31:0] _cp0_io_exception_type_i; // @[myCPU.scala 123:22]
  wire  _cp0_io_in_delayslot; // @[myCPU.scala 123:22]
  wire [1:0] _cp0_io_in_branchjump_jr; // @[myCPU.scala 123:22]
  wire [31:0] _cp0_io_return_pc; // @[myCPU.scala 123:22]
  wire  _cp0_io_exception; // @[myCPU.scala 123:22]
  wire [31:0] _cp0_io_cp0_read_data; // @[myCPU.scala 123:22]
  wire [31:0] _cp0_io_epc; // @[myCPU.scala 123:22]
  wire [5:0] _cp0_io_cp0_status; // @[myCPU.scala 123:22]
  wire  _cp0_io_Int_able; // @[myCPU.scala 123:22]
  wire [7:0] _cp0_io_asid; // @[myCPU.scala 123:22]
  wire [18:0] _cp0_io_cp0_tlb_read_data_vaddr; // @[myCPU.scala 123:22]
  wire [7:0] _cp0_io_cp0_tlb_read_data_asid; // @[myCPU.scala 123:22]
  wire  _cp0_io_cp0_tlb_read_data_g; // @[myCPU.scala 123:22]
  wire [19:0] _cp0_io_cp0_tlb_read_data_paddr_0; // @[myCPU.scala 123:22]
  wire [19:0] _cp0_io_cp0_tlb_read_data_paddr_1; // @[myCPU.scala 123:22]
  wire [2:0] _cp0_io_cp0_tlb_read_data_c_0; // @[myCPU.scala 123:22]
  wire [2:0] _cp0_io_cp0_tlb_read_data_c_1; // @[myCPU.scala 123:22]
  wire  _cp0_io_cp0_tlb_read_data_d_0; // @[myCPU.scala 123:22]
  wire  _cp0_io_cp0_tlb_read_data_d_1; // @[myCPU.scala 123:22]
  wire  _cp0_io_cp0_tlb_read_data_v_0; // @[myCPU.scala 123:22]
  wire  _cp0_io_cp0_tlb_read_data_v_1; // @[myCPU.scala 123:22]
  wire [18:0] _cp0_io_cp0_tlb_write_data_vaddr; // @[myCPU.scala 123:22]
  wire [7:0] _cp0_io_cp0_tlb_write_data_asid; // @[myCPU.scala 123:22]
  wire  _cp0_io_cp0_tlb_write_data_g; // @[myCPU.scala 123:22]
  wire [19:0] _cp0_io_cp0_tlb_write_data_paddr_0; // @[myCPU.scala 123:22]
  wire [19:0] _cp0_io_cp0_tlb_write_data_paddr_1; // @[myCPU.scala 123:22]
  wire [2:0] _cp0_io_cp0_tlb_write_data_c_0; // @[myCPU.scala 123:22]
  wire [2:0] _cp0_io_cp0_tlb_write_data_c_1; // @[myCPU.scala 123:22]
  wire  _cp0_io_cp0_tlb_write_data_d_0; // @[myCPU.scala 123:22]
  wire  _cp0_io_cp0_tlb_write_data_d_1; // @[myCPU.scala 123:22]
  wire  _cp0_io_cp0_tlb_write_data_v_0; // @[myCPU.scala 123:22]
  wire  _cp0_io_cp0_tlb_write_data_v_1; // @[myCPU.scala 123:22]
  wire  _cp0_io_cp0_tlb_write_en; // @[myCPU.scala 123:22]
  wire  _cp0_io_cp0_index_tlb_write_able; // @[myCPU.scala 123:22]
  wire  _cu_reset; // @[myCPU.scala 124:22]
  wire [31:0] _cu_io1_InstrD; // @[myCPU.scala 124:22]
  wire  _cu_io1_BadInstrD; // @[myCPU.scala 124:22]
  wire  _cu_io1_BreakD; // @[myCPU.scala 124:22]
  wire  _cu_io1_SysCallD; // @[myCPU.scala 124:22]
  wire  _cu_io1_EretD; // @[myCPU.scala 124:22]
  wire [2:0] _cu_io1_Tlb_Control; // @[myCPU.scala 124:22]
  wire  _cu_io1_commit_cache_ins; // @[myCPU.scala 124:22]
  wire  _cu_io1_dmem_addr_cal; // @[myCPU.scala 124:22]
  wire  _cu_io_RegWriteD; // @[myCPU.scala 124:22]
  wire  _cu_io_MemToRegD; // @[myCPU.scala 124:22]
  wire  _cu_io_MemWriteD; // @[myCPU.scala 124:22]
  wire [23:0] _cu_io_ALUCtrlD; // @[myCPU.scala 124:22]
  wire [1:0] _cu_io_ALUSrcD; // @[myCPU.scala 124:22]
  wire [1:0] _cu_io_RegDstD; // @[myCPU.scala 124:22]
  wire  _cu_io_ImmUnsigned; // @[myCPU.scala 124:22]
  wire  _cu_io_LinkD; // @[myCPU.scala 124:22]
  wire [1:0] _cu_io_HiLoWriteD; // @[myCPU.scala 124:22]
  wire [1:0] _cu_io_HiLoToRegD; // @[myCPU.scala 124:22]
  wire  _cu_io_CP0WriteD; // @[myCPU.scala 124:22]
  wire  _cu_io_CP0ToRegD; // @[myCPU.scala 124:22]
  wire  _cu_io_LoadUnsignedD; // @[myCPU.scala 124:22]
  wire [1:0] _cu_io_MemWidthD; // @[myCPU.scala 124:22]
  wire [1:0] _cu_io_MemRLD; // @[myCPU.scala 124:22]
  wire  _dmem_io_data_ok; // @[myCPU.scala 125:23]
  wire [31:0] _dmem_io_rdata; // @[myCPU.scala 125:23]
  wire [31:0] _dmem_io_Physisc_Address; // @[myCPU.scala 125:23]
  wire [1:0] _dmem_io_WIDTH; // @[myCPU.scala 125:23]
  wire  _dmem_io_SIGN; // @[myCPU.scala 125:23]
  wire [31:0] _dmem_io_RD; // @[myCPU.scala 125:23]
  wire  _dmem_io_data_pending; // @[myCPU.scala 125:23]
  wire  _dmemreq_io_en; // @[myCPU.scala 126:26]
  wire  _dmemreq_io_MemWriteE; // @[myCPU.scala 126:26]
  wire  _dmemreq_io_MemToRegE; // @[myCPU.scala 126:26]
  wire [1:0] _dmemreq_io_MemWidthE; // @[myCPU.scala 126:26]
  wire [31:0] _dmemreq_io_VAddrE; // @[myCPU.scala 126:26]
  wire [31:0] _dmemreq_io_WriteDataE; // @[myCPU.scala 126:26]
  wire [1:0] _dmemreq_io_memrl; // @[myCPU.scala 126:26]
  wire  _dmemreq_io_req; // @[myCPU.scala 126:26]
  wire  _dmemreq_io_wr; // @[myCPU.scala 126:26]
  wire [1:0] _dmemreq_io_size; // @[myCPU.scala 126:26]
  wire [31:0] _dmemreq_io_addr; // @[myCPU.scala 126:26]
  wire [31:0] _dmemreq_io_wdata; // @[myCPU.scala 126:26]
  wire [3:0] _dmemreq_io_wstrb; // @[myCPU.scala 126:26]
  wire  _ex2mem_clock; // @[myCPU.scala 127:26]
  wire  _ex2mem_reset; // @[myCPU.scala 127:26]
  wire  _ex2mem_io1_RegWriteE; // @[myCPU.scala 127:26]
  wire  _ex2mem_io1_MemToRegE; // @[myCPU.scala 127:26]
  wire  _ex2mem_io1_LoadUnsignedE; // @[myCPU.scala 127:26]
  wire [1:0] _ex2mem_io1_MemWidthE; // @[myCPU.scala 127:26]
  wire [1:0] _ex2mem_io1_HiLoWriteE; // @[myCPU.scala 127:26]
  wire  _ex2mem_io1_CP0WriteE; // @[myCPU.scala 127:26]
  wire [4:0] _ex2mem_io1_WriteCP0AddrE; // @[myCPU.scala 127:26]
  wire [2:0] _ex2mem_io1_WriteCP0SelE; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io1_PCE; // @[myCPU.scala 127:26]
  wire  _ex2mem_io1_InDelaySlotE; // @[myCPU.scala 127:26]
  wire [1:0] _ex2mem_io1_MemRLE; // @[myCPU.scala 127:26]
  wire [1:0] _ex2mem_io1_BranchJump_JrE; // @[myCPU.scala 127:26]
  wire [2:0] _ex2mem_io1_Tlb_Control; // @[myCPU.scala 127:26]
  wire  _ex2mem_io_en; // @[myCPU.scala 127:26]
  wire  _ex2mem_io_clr; // @[myCPU.scala 127:26]
  wire [4:0] _ex2mem_io_WriteRegE; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_PhyAddrE; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_HiLoOutE; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_HiInE; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_LoInE; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_WriteCP0HiLoDataE; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_BadVAddrE; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_ExceptionTypeE; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_RtE; // @[myCPU.scala 127:26]
  wire  _ex2mem_io_RegWriteM; // @[myCPU.scala 127:26]
  wire  _ex2mem_io_MemToRegM; // @[myCPU.scala 127:26]
  wire [4:0] _ex2mem_io_WriteRegM; // @[myCPU.scala 127:26]
  wire  _ex2mem_io_LoadUnsignedM; // @[myCPU.scala 127:26]
  wire [1:0] _ex2mem_io_MemWidthM; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_PhyAddrM; // @[myCPU.scala 127:26]
  wire [1:0] _ex2mem_io_HiLoWriteM; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_HiLoOutM; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_HiInM; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_LoInM; // @[myCPU.scala 127:26]
  wire  _ex2mem_io_CP0WriteM; // @[myCPU.scala 127:26]
  wire [4:0] _ex2mem_io_WriteCP0AddrM; // @[myCPU.scala 127:26]
  wire [2:0] _ex2mem_io_WriteCP0SelM; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_WriteCP0HiLoDataM; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_PCM; // @[myCPU.scala 127:26]
  wire  _ex2mem_io_InDelaySlotM; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_BadVAddrM; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_ExceptionTypeM_Out; // @[myCPU.scala 127:26]
  wire [1:0] _ex2mem_io_MemRLM; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_RtM; // @[myCPU.scala 127:26]
  wire [1:0] _ex2mem_io_BranchJump_JrM; // @[myCPU.scala 127:26]
  wire [2:0] _ex2mem_io_Tlb_ControlM; // @[myCPU.scala 127:26]
  wire  _mem2mem2_clock; // @[myCPU.scala 128:28]
  wire  _mem2mem2_reset; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io1_RegWriteE; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io1_MemToRegE; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io1_LoadUnsignedE; // @[myCPU.scala 128:28]
  wire [1:0] _mem2mem2_io1_MemWidthE; // @[myCPU.scala 128:28]
  wire [1:0] _mem2mem2_io1_HiLoWriteE; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io1_CP0WriteE; // @[myCPU.scala 128:28]
  wire [4:0] _mem2mem2_io1_WriteCP0AddrE; // @[myCPU.scala 128:28]
  wire [2:0] _mem2mem2_io1_WriteCP0SelE; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io1_PCE; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io1_InDelaySlotE; // @[myCPU.scala 128:28]
  wire [1:0] _mem2mem2_io1_MemRLE; // @[myCPU.scala 128:28]
  wire [1:0] _mem2mem2_io1_BranchJump_JrE; // @[myCPU.scala 128:28]
  wire [2:0] _mem2mem2_io1_Tlb_Control; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io_en; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io_clr; // @[myCPU.scala 128:28]
  wire [4:0] _mem2mem2_io_WriteRegE; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_PhyAddrE; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_HiLoOutE; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_HiInE; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_LoInE; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_WriteCP0HiLoDataE; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_BadVAddrE; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_ExceptionTypeE; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_RtE; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io_RegWriteM; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io_MemToRegM; // @[myCPU.scala 128:28]
  wire [4:0] _mem2mem2_io_WriteRegM; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io_LoadUnsignedM; // @[myCPU.scala 128:28]
  wire [1:0] _mem2mem2_io_MemWidthM; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_PhyAddrM; // @[myCPU.scala 128:28]
  wire [1:0] _mem2mem2_io_HiLoWriteM; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_HiLoOutM; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_HiInM; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_LoInM; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io_CP0WriteM; // @[myCPU.scala 128:28]
  wire [4:0] _mem2mem2_io_WriteCP0AddrM; // @[myCPU.scala 128:28]
  wire [2:0] _mem2mem2_io_WriteCP0SelM; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_WriteCP0HiLoDataM; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_PCM; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io_InDelaySlotM; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_BadVAddrM; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_ExceptionTypeM_Out; // @[myCPU.scala 128:28]
  wire [1:0] _mem2mem2_io_MemRLM; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_RtM; // @[myCPU.scala 128:28]
  wire [1:0] _mem2mem2_io_BranchJump_JrM; // @[myCPU.scala 128:28]
  wire [2:0] _mem2mem2_io_Tlb_ControlM; // @[myCPU.scala 128:28]
  wire  _hilo_clock; // @[myCPU.scala 129:26]
  wire  _hilo_reset; // @[myCPU.scala 129:26]
  wire [1:0] _hilo_io_we; // @[myCPU.scala 129:26]
  wire [31:0] _hilo_io_hi_i; // @[myCPU.scala 129:26]
  wire [31:0] _hilo_io_lo_i; // @[myCPU.scala 129:26]
  wire [31:0] _hilo_io_hi_o; // @[myCPU.scala 129:26]
  wire [31:0] _hilo_io_lo_o; // @[myCPU.scala 129:26]
  wire  _id2ex_clock; // @[myCPU.scala 130:26]
  wire  _id2ex_reset; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_RegWriteD; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_MemToRegD; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_MemWriteD; // @[myCPU.scala 130:26]
  wire [23:0] _id2ex_io1_ALUCtrlD; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io1_ALUSrcD; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io1_RegDstD; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_LinkD; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io1_HiLoWriteD; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io1_HiLoToRegD; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_CP0WriteD; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_CP0ToRegD; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_LoadUnsignedD; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io1_MemWidthD; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io1_MemRLD; // @[myCPU.scala 130:26]
  wire  _id2ex_io2_RegWriteE; // @[myCPU.scala 130:26]
  wire  _id2ex_io2_MemToRegE; // @[myCPU.scala 130:26]
  wire  _id2ex_io2_MemWriteE; // @[myCPU.scala 130:26]
  wire [23:0] _id2ex_io2_ALUCtrlE; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io2_ALUSrcE; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io2_RegDstE; // @[myCPU.scala 130:26]
  wire  _id2ex_io2_LinkE; // @[myCPU.scala 130:26]
  wire [31:0] _id2ex_io2_PCPlus8E; // @[myCPU.scala 130:26]
  wire  _id2ex_io2_LoadUnsignedE; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io2_MemWidthE; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io2_HiLoWriteE; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io2_HiLoToRegE; // @[myCPU.scala 130:26]
  wire  _id2ex_io2_CP0WriteE; // @[myCPU.scala 130:26]
  wire [4:0] _id2ex_io2_WriteCP0AddrE; // @[myCPU.scala 130:26]
  wire [2:0] _id2ex_io2_WriteCP0SelE; // @[myCPU.scala 130:26]
  wire [4:0] _id2ex_io2_ReadCP0AddrE; // @[myCPU.scala 130:26]
  wire [2:0] _id2ex_io2_ReadCP0SelE; // @[myCPU.scala 130:26]
  wire [31:0] _id2ex_io2_PCE; // @[myCPU.scala 130:26]
  wire  _id2ex_io2_InDelaySlotE; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io2_MemRLE; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io2_BranchJump_JrE; // @[myCPU.scala 130:26]
  wire [2:0] _id2ex_io2_Tlb_Control; // @[myCPU.scala 130:26]
  wire  _id2ex_io_en; // @[myCPU.scala 130:26]
  wire  _id2ex_io_clr; // @[myCPU.scala 130:26]
  wire  _id2ex_io_CP0ToRegE_Out; // @[myCPU.scala 130:26]
  wire [31:0] _id2ex_io_RD1D; // @[myCPU.scala 130:26]
  wire [31:0] _id2ex_io_RD2D; // @[myCPU.scala 130:26]
  wire [4:0] _id2ex_io_RsD; // @[myCPU.scala 130:26]
  wire [4:0] _id2ex_io_RtD; // @[myCPU.scala 130:26]
  wire [4:0] _id2ex_io_RdD; // @[myCPU.scala 130:26]
  wire [31:0] _id2ex_io_ImmD; // @[myCPU.scala 130:26]
  wire [31:0] _id2ex_io_PCPlus8D; // @[myCPU.scala 130:26]
  wire [4:0] _id2ex_io_WriteCP0AddrD; // @[myCPU.scala 130:26]
  wire [2:0] _id2ex_io_WriteCP0SelD; // @[myCPU.scala 130:26]
  wire [4:0] _id2ex_io_ReadCP0AddrD; // @[myCPU.scala 130:26]
  wire [2:0] _id2ex_io_ReadCP0SelD; // @[myCPU.scala 130:26]
  wire [31:0] _id2ex_io_PCD; // @[myCPU.scala 130:26]
  wire  _id2ex_io_InDelaySlotD; // @[myCPU.scala 130:26]
  wire [31:0] _id2ex_io_ExceptionTypeD; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io_BranchJump_JrD; // @[myCPU.scala 130:26]
  wire [31:0] _id2ex_io_BadVaddrD; // @[myCPU.scala 130:26]
  wire [2:0] _id2ex_io_Tlb_Control; // @[myCPU.scala 130:26]
  wire [31:0] _id2ex_io_RD1E; // @[myCPU.scala 130:26]
  wire [31:0] _id2ex_io_RD2E; // @[myCPU.scala 130:26]
  wire [4:0] _id2ex_io_RsE; // @[myCPU.scala 130:26]
  wire [4:0] _id2ex_io_RtE; // @[myCPU.scala 130:26]
  wire [4:0] _id2ex_io_RdE; // @[myCPU.scala 130:26]
  wire [31:0] _id2ex_io_ImmE; // @[myCPU.scala 130:26]
  wire [31:0] _id2ex_io_BadVaddrE; // @[myCPU.scala 130:26]
  wire [31:0] _id2ex_io_ExceptionTypeE_Out; // @[myCPU.scala 130:26]
  wire  _if2id_clock; // @[myCPU.scala 131:26]
  wire  _if2id_reset; // @[myCPU.scala 131:26]
  wire  _if2id_io_en; // @[myCPU.scala 131:26]
  wire  _if2id_io_clr; // @[myCPU.scala 131:26]
  wire [31:0] _if2id_io_InstrF; // @[myCPU.scala 131:26]
  wire [31:0] _if2id_io_PCPlus4F; // @[myCPU.scala 131:26]
  wire [31:0] _if2id_io_PCPlus8F; // @[myCPU.scala 131:26]
  wire [31:0] _if2id_io_PCF; // @[myCPU.scala 131:26]
  wire [1:0] _if2id_io_ExceptionTypeF; // @[myCPU.scala 131:26]
  wire  _if2id_io_NextDelaySlotD; // @[myCPU.scala 131:26]
  wire [31:0] _if2id_io_InstrD; // @[myCPU.scala 131:26]
  wire [31:0] _if2id_io_PCPlus4D; // @[myCPU.scala 131:26]
  wire [31:0] _if2id_io_PCPlus8D; // @[myCPU.scala 131:26]
  wire  _if2id_io_InDelaySlotD; // @[myCPU.scala 131:26]
  wire [31:0] _if2id_io_PCD; // @[myCPU.scala 131:26]
  wire [1:0] _if2id_io_ExceptionTypeD_Out; // @[myCPU.scala 131:26]
  wire  _mem22wb_clock; // @[myCPU.scala 133:27]
  wire  _mem22wb_reset; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_en; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_clr; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_RegWriteM; // @[myCPU.scala 133:27]
  wire [31:0] _mem22wb_io_ResultM; // @[myCPU.scala 133:27]
  wire [4:0] _mem22wb_io_WriteRegM; // @[myCPU.scala 133:27]
  wire [1:0] _mem22wb_io_HiLoWriteM; // @[myCPU.scala 133:27]
  wire [31:0] _mem22wb_io_HiInM; // @[myCPU.scala 133:27]
  wire [31:0] _mem22wb_io_LoInM; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_CP0WriteM; // @[myCPU.scala 133:27]
  wire [4:0] _mem22wb_io_WriteCP0AddrM; // @[myCPU.scala 133:27]
  wire [2:0] _mem22wb_io_WriteCP0SelM; // @[myCPU.scala 133:27]
  wire [31:0] _mem22wb_io_WriteCP0HiLoDataM; // @[myCPU.scala 133:27]
  wire [31:0] _mem22wb_io_PCM; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_InDelaySlotM; // @[myCPU.scala 133:27]
  wire [31:0] _mem22wb_io_BadVAddrM; // @[myCPU.scala 133:27]
  wire [31:0] _mem22wb_io_ExceptionTypeM; // @[myCPU.scala 133:27]
  wire [1:0] _mem22wb_io_BranchJump_JrM; // @[myCPU.scala 133:27]
  wire [2:0] _mem22wb_io_Tlb_ControlM; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_RegWriteW_Out; // @[myCPU.scala 133:27]
  wire [31:0] _mem22wb_io_ResultW; // @[myCPU.scala 133:27]
  wire [4:0] _mem22wb_io_WriteRegW; // @[myCPU.scala 133:27]
  wire [1:0] _mem22wb_io_HiLoWriteW; // @[myCPU.scala 133:27]
  wire [31:0] _mem22wb_io_HiInW; // @[myCPU.scala 133:27]
  wire [31:0] _mem22wb_io_LoInW; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_CP0WriteW; // @[myCPU.scala 133:27]
  wire [4:0] _mem22wb_io_WriteCP0AddrW; // @[myCPU.scala 133:27]
  wire [2:0] _mem22wb_io_WriteCP0SelW; // @[myCPU.scala 133:27]
  wire [31:0] _mem22wb_io_WriteCP0HiLoDataW; // @[myCPU.scala 133:27]
  wire [31:0] _mem22wb_io_PCW; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_InDelaySlotW; // @[myCPU.scala 133:27]
  wire [31:0] _mem22wb_io_BadVAddrW; // @[myCPU.scala 133:27]
  wire [31:0] _mem22wb_io_ExceptionTypeW_Out; // @[myCPU.scala 133:27]
  wire [1:0] _mem22wb_io_BranchJump_JrW; // @[myCPU.scala 133:27]
  wire [2:0] _mem22wb_io_Tlb_ControlW; // @[myCPU.scala 133:27]
  wire [31:0] _addr_cal_io_d_vaddr; // @[myCPU.scala 134:31]
  wire [1:0] _addr_cal_io_d_width; // @[myCPU.scala 134:31]
  wire [1:0] _addr_cal_io_d_memrl; // @[myCPU.scala 134:31]
  wire [31:0] _addr_cal_io_d_paddr; // @[myCPU.scala 134:31]
  wire  _addr_cal_io_d_cached; // @[myCPU.scala 134:31]
  wire  _addr_cal_io_d_unaligned; // @[myCPU.scala 134:31]
  wire  _muldiv_clock; // @[myCPU.scala 135:26]
  wire  _muldiv_reset; // @[myCPU.scala 135:26]
  wire  _muldiv_io_en; // @[myCPU.scala 135:26]
  wire [4:0] _muldiv_io_ctrl; // @[myCPU.scala 135:26]
  wire [31:0] _muldiv_io_in1; // @[myCPU.scala 135:26]
  wire [31:0] _muldiv_io_in2; // @[myCPU.scala 135:26]
  wire [31:0] _muldiv_io_hi; // @[myCPU.scala 135:26]
  wire [31:0] _muldiv_io_lo; // @[myCPU.scala 135:26]
  wire  _muldiv_io_pending; // @[myCPU.scala 135:26]
  wire  _regfile_clock; // @[myCPU.scala 137:26]
  wire  _regfile_reset; // @[myCPU.scala 137:26]
  wire [4:0] _regfile_io_A1; // @[myCPU.scala 137:26]
  wire [4:0] _regfile_io_A2; // @[myCPU.scala 137:26]
  wire  _regfile_io_WE3; // @[myCPU.scala 137:26]
  wire [4:0] _regfile_io_A3; // @[myCPU.scala 137:26]
  wire [31:0] _regfile_io_WD3; // @[myCPU.scala 137:26]
  wire [31:0] _regfile_io_RD1; // @[myCPU.scala 137:26]
  wire [31:0] _regfile_io_RD2; // @[myCPU.scala 137:26]
  wire  fifo_clock; // @[myCPU.scala 139:29]
  wire  fifo_reset; // @[myCPU.scala 139:29]
  wire [1:0] fifo_io_read_en; // @[myCPU.scala 139:29]
  wire [1:0] fifo_io_write_en; // @[myCPU.scala 139:29]
  wire [135:0] fifo_io_read_out_0; // @[myCPU.scala 139:29]
  wire [135:0] fifo_io_write_in_0; // @[myCPU.scala 139:29]
  wire  fifo_io_full; // @[myCPU.scala 139:29]
  wire  fifo_io_empty; // @[myCPU.scala 139:29]
  wire  fifo_io_point_write_en; // @[myCPU.scala 139:29]
  wire  fifo_io_point_flush; // @[myCPU.scala 139:29]
  wire  stage_fec_1_pc_L_clock; // @[myCPU.scala 403:34]
  wire  stage_fec_1_pc_L_reset; // @[myCPU.scala 403:34]
  wire  stage_fec_1_pc_L_io_stall; // @[myCPU.scala 403:34]
  wire  stage_fec_1_pc_L_io_flush; // @[myCPU.scala 403:34]
  wire [31:0] stage_fec_1_pc_L_io_in_pc_value_in; // @[myCPU.scala 403:34]
  wire [31:0] stage_fec_1_pc_L_io_out_pc_value_out; // @[myCPU.scala 403:34]
  wire  stage_fec_1_pc_M_clock; // @[myCPU.scala 404:34]
  wire  stage_fec_1_pc_M_reset; // @[myCPU.scala 404:34]
  wire  stage_fec_1_pc_M_io_stall; // @[myCPU.scala 404:34]
  wire  stage_fec_1_pc_M_io_flush; // @[myCPU.scala 404:34]
  wire [31:0] stage_fec_1_pc_M_io_in_pc_value_in; // @[myCPU.scala 404:34]
  wire [31:0] stage_fec_1_pc_M_io_out_pc_value_out; // @[myCPU.scala 404:34]
  wire  stage_fec_1_pc_R_clock; // @[myCPU.scala 405:34]
  wire  stage_fec_1_pc_R_reset; // @[myCPU.scala 405:34]
  wire  stage_fec_1_pc_R_io_stall; // @[myCPU.scala 405:34]
  wire  stage_fec_1_pc_R_io_flush; // @[myCPU.scala 405:34]
  wire [31:0] stage_fec_1_pc_R_io_in_pc_value_in; // @[myCPU.scala 405:34]
  wire [31:0] stage_fec_1_pc_R_io_out_pc_value_out; // @[myCPU.scala 405:34]
  wire  branch_prediction_with_blockram_clock; // @[myCPU.scala 434:21]
  wire  branch_prediction_with_blockram_reset; // @[myCPU.scala 434:21]
  wire [31:0] branch_prediction_with_blockram_io_pc; // @[myCPU.scala 434:21]
  wire [31:0] branch_prediction_with_blockram_io_write_pc; // @[myCPU.scala 434:21]
  wire [3:0] branch_prediction_with_blockram_io_aw_pht_ways_addr; // @[myCPU.scala 434:21]
  wire [6:0] branch_prediction_with_blockram_io_aw_pht_addr; // @[myCPU.scala 434:21]
  wire [6:0] branch_prediction_with_blockram_io_aw_bht_addr; // @[myCPU.scala 434:21]
  wire [31:0] branch_prediction_with_blockram_io_aw_target_addr; // @[myCPU.scala 434:21]
  wire  branch_prediction_with_blockram_io_btb_write; // @[myCPU.scala 434:21]
  wire  branch_prediction_with_blockram_io_bht_write; // @[myCPU.scala 434:21]
  wire  branch_prediction_with_blockram_io_pht_write; // @[myCPU.scala 434:21]
  wire [6:0] branch_prediction_with_blockram_io_bht_in; // @[myCPU.scala 434:21]
  wire [7:0] branch_prediction_with_blockram_io_pht_in; // @[myCPU.scala 434:21]
  wire [1:0] branch_prediction_with_blockram_io_out_L; // @[myCPU.scala 434:21]
  wire  branch_prediction_with_blockram_io_pre_L; // @[myCPU.scala 434:21]
  wire [6:0] branch_prediction_with_blockram_io_bht_L; // @[myCPU.scala 434:21]
  wire  branch_prediction_with_blockram_io_btb_hit_0; // @[myCPU.scala 434:21]
  wire [31:0] branch_prediction_with_blockram_io_pre_target_L; // @[myCPU.scala 434:21]
  wire  branch_prediction_with_blockram_io_stage2_stall; // @[myCPU.scala 434:21]
  wire  branch_prediction_with_blockram_io_stage2_flush; // @[myCPU.scala 434:21]
  wire [7:0] branch_prediction_with_blockram_io_pht_out; // @[myCPU.scala 434:21]
  wire [6:0] branch_prediction_with_blockram_io_lookup_data_0; // @[myCPU.scala 434:21]
  wire  stage_fec_2_pc_L_clock; // @[myCPU.scala 503:34]
  wire  stage_fec_2_pc_L_reset; // @[myCPU.scala 503:34]
  wire  stage_fec_2_pc_L_io_stall; // @[myCPU.scala 503:34]
  wire  stage_fec_2_pc_L_io_flush; // @[myCPU.scala 503:34]
  wire [31:0] stage_fec_2_pc_L_io_in_pc_value_in; // @[myCPU.scala 503:34]
  wire [31:0] stage_fec_2_pc_L_io_out_pc_value_out; // @[myCPU.scala 503:34]
  wire  stage_fec_2_pc_M_clock; // @[myCPU.scala 504:34]
  wire  stage_fec_2_pc_M_reset; // @[myCPU.scala 504:34]
  wire  stage_fec_2_pc_M_io_stall; // @[myCPU.scala 504:34]
  wire  stage_fec_2_pc_M_io_flush; // @[myCPU.scala 504:34]
  wire [31:0] stage_fec_2_pc_M_io_in_pc_value_in; // @[myCPU.scala 504:34]
  wire [31:0] stage_fec_2_pc_M_io_out_pc_value_out; // @[myCPU.scala 504:34]
  wire  stage_fec_2_pc_R_clock; // @[myCPU.scala 505:34]
  wire  stage_fec_2_pc_R_reset; // @[myCPU.scala 505:34]
  wire  stage_fec_2_pc_R_io_stall; // @[myCPU.scala 505:34]
  wire  stage_fec_2_pc_R_io_flush; // @[myCPU.scala 505:34]
  wire [31:0] stage_fec_2_pc_R_io_in_pc_value_in; // @[myCPU.scala 505:34]
  wire [31:0] stage_fec_2_pc_R_io_out_pc_value_out; // @[myCPU.scala 505:34]
  wire  id_bru_state_clock; // @[myCPU.scala 652:27]
  wire  id_bru_state_reset; // @[myCPU.scala 652:27]
  wire  id_bru_state_io_stall; // @[myCPU.scala 652:27]
  wire  id_bru_state_io_flush; // @[myCPU.scala 652:27]
  wire [1:0] id_bru_state_io_in_pht; // @[myCPU.scala 652:27]
  wire [6:0] id_bru_state_io_in_bht; // @[myCPU.scala 652:27]
  wire [3:0] id_bru_state_io_in_hashcode; // @[myCPU.scala 652:27]
  wire [31:0] id_bru_state_io_in_target_pc; // @[myCPU.scala 652:27]
  wire [6:0] id_bru_state_io_in_lookup_data; // @[myCPU.scala 652:27]
  wire [7:0] id_bru_state_io_in_pht_lookup_value; // @[myCPU.scala 652:27]
  wire [1:0] id_bru_state_io_out_pht; // @[myCPU.scala 652:27]
  wire [6:0] id_bru_state_io_out_bht; // @[myCPU.scala 652:27]
  wire [3:0] id_bru_state_io_out_hashcode; // @[myCPU.scala 652:27]
  wire [31:0] id_bru_state_io_out_target_pc; // @[myCPU.scala 652:27]
  wire [6:0] id_bru_state_io_out_lookup_data; // @[myCPU.scala 652:27]
  wire [7:0] id_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 652:27]
  wire  ex_bru_state_clock; // @[myCPU.scala 656:27]
  wire  ex_bru_state_reset; // @[myCPU.scala 656:27]
  wire  ex_bru_state_io_stall; // @[myCPU.scala 656:27]
  wire  ex_bru_state_io_flush; // @[myCPU.scala 656:27]
  wire [1:0] ex_bru_state_io_in_pht; // @[myCPU.scala 656:27]
  wire [6:0] ex_bru_state_io_in_bht; // @[myCPU.scala 656:27]
  wire [3:0] ex_bru_state_io_in_hashcode; // @[myCPU.scala 656:27]
  wire [31:0] ex_bru_state_io_in_target_pc; // @[myCPU.scala 656:27]
  wire [6:0] ex_bru_state_io_in_lookup_data; // @[myCPU.scala 656:27]
  wire [7:0] ex_bru_state_io_in_pht_lookup_value; // @[myCPU.scala 656:27]
  wire [1:0] ex_bru_state_io_out_pht; // @[myCPU.scala 656:27]
  wire [6:0] ex_bru_state_io_out_bht; // @[myCPU.scala 656:27]
  wire [3:0] ex_bru_state_io_out_hashcode; // @[myCPU.scala 656:27]
  wire [31:0] ex_bru_state_io_out_target_pc; // @[myCPU.scala 656:27]
  wire [6:0] ex_bru_state_io_out_lookup_data; // @[myCPU.scala 656:27]
  wire [7:0] ex_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 656:27]
  wire  mem_bru_state_clock; // @[myCPU.scala 660:28]
  wire  mem_bru_state_reset; // @[myCPU.scala 660:28]
  wire  mem_bru_state_io_stall; // @[myCPU.scala 660:28]
  wire  mem_bru_state_io_flush; // @[myCPU.scala 660:28]
  wire [1:0] mem_bru_state_io_in_pht; // @[myCPU.scala 660:28]
  wire [6:0] mem_bru_state_io_in_bht; // @[myCPU.scala 660:28]
  wire [3:0] mem_bru_state_io_in_hashcode; // @[myCPU.scala 660:28]
  wire [31:0] mem_bru_state_io_in_target_pc; // @[myCPU.scala 660:28]
  wire [6:0] mem_bru_state_io_in_lookup_data; // @[myCPU.scala 660:28]
  wire [7:0] mem_bru_state_io_in_pht_lookup_value; // @[myCPU.scala 660:28]
  wire [1:0] mem_bru_state_io_out_pht; // @[myCPU.scala 660:28]
  wire [6:0] mem_bru_state_io_out_bht; // @[myCPU.scala 660:28]
  wire [3:0] mem_bru_state_io_out_hashcode; // @[myCPU.scala 660:28]
  wire [31:0] mem_bru_state_io_out_target_pc; // @[myCPU.scala 660:28]
  wire [6:0] mem_bru_state_io_out_lookup_data; // @[myCPU.scala 660:28]
  wire [7:0] mem_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 660:28]
  wire  mem2_bru_state_clock; // @[myCPU.scala 664:29]
  wire  mem2_bru_state_reset; // @[myCPU.scala 664:29]
  wire  mem2_bru_state_io_stall; // @[myCPU.scala 664:29]
  wire  mem2_bru_state_io_flush; // @[myCPU.scala 664:29]
  wire [1:0] mem2_bru_state_io_in_pht; // @[myCPU.scala 664:29]
  wire [6:0] mem2_bru_state_io_in_bht; // @[myCPU.scala 664:29]
  wire [3:0] mem2_bru_state_io_in_hashcode; // @[myCPU.scala 664:29]
  wire [31:0] mem2_bru_state_io_in_target_pc; // @[myCPU.scala 664:29]
  wire [6:0] mem2_bru_state_io_in_lookup_data; // @[myCPU.scala 664:29]
  wire [7:0] mem2_bru_state_io_in_pht_lookup_value; // @[myCPU.scala 664:29]
  wire [1:0] mem2_bru_state_io_out_pht; // @[myCPU.scala 664:29]
  wire [6:0] mem2_bru_state_io_out_bht; // @[myCPU.scala 664:29]
  wire [3:0] mem2_bru_state_io_out_hashcode; // @[myCPU.scala 664:29]
  wire [31:0] mem2_bru_state_io_out_target_pc; // @[myCPU.scala 664:29]
  wire [6:0] mem2_bru_state_io_out_lookup_data; // @[myCPU.scala 664:29]
  wire [7:0] mem2_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 664:29]
  wire  wb_bru_state_clock; // @[myCPU.scala 668:27]
  wire  wb_bru_state_reset; // @[myCPU.scala 668:27]
  wire  wb_bru_state_io_stall; // @[myCPU.scala 668:27]
  wire  wb_bru_state_io_flush; // @[myCPU.scala 668:27]
  wire [1:0] wb_bru_state_io_in_pht; // @[myCPU.scala 668:27]
  wire [6:0] wb_bru_state_io_in_bht; // @[myCPU.scala 668:27]
  wire [3:0] wb_bru_state_io_in_hashcode; // @[myCPU.scala 668:27]
  wire [31:0] wb_bru_state_io_in_target_pc; // @[myCPU.scala 668:27]
  wire [6:0] wb_bru_state_io_in_lookup_data; // @[myCPU.scala 668:27]
  wire [7:0] wb_bru_state_io_in_pht_lookup_value; // @[myCPU.scala 668:27]
  wire [1:0] wb_bru_state_io_out_pht; // @[myCPU.scala 668:27]
  wire [6:0] wb_bru_state_io_out_bht; // @[myCPU.scala 668:27]
  wire [3:0] wb_bru_state_io_out_hashcode; // @[myCPU.scala 668:27]
  wire [31:0] wb_bru_state_io_out_target_pc; // @[myCPU.scala 668:27]
  wire [6:0] wb_bru_state_io_out_lookup_data; // @[myCPU.scala 668:27]
  wire [7:0] wb_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 668:27]
  wire  tlb_data_register_clock; // @[myCPU.scala 971:30]
  wire  tlb_data_register_reset; // @[myCPU.scala 971:30]
  wire  tlb_data_register_io_flush; // @[myCPU.scala 971:30]
  wire  tlb_data_register_io_stall; // @[myCPU.scala 971:30]
  wire [18:0] tlb_data_register_io_tlb_read_data_vaddr; // @[myCPU.scala 971:30]
  wire [7:0] tlb_data_register_io_tlb_read_data_asid; // @[myCPU.scala 971:30]
  wire  tlb_data_register_io_tlb_read_data_g; // @[myCPU.scala 971:30]
  wire [19:0] tlb_data_register_io_tlb_read_data_paddr_0; // @[myCPU.scala 971:30]
  wire [19:0] tlb_data_register_io_tlb_read_data_paddr_1; // @[myCPU.scala 971:30]
  wire [2:0] tlb_data_register_io_tlb_read_data_c_0; // @[myCPU.scala 971:30]
  wire [2:0] tlb_data_register_io_tlb_read_data_c_1; // @[myCPU.scala 971:30]
  wire  tlb_data_register_io_tlb_read_data_d_0; // @[myCPU.scala 971:30]
  wire  tlb_data_register_io_tlb_read_data_d_1; // @[myCPU.scala 971:30]
  wire  tlb_data_register_io_tlb_read_data_v_0; // @[myCPU.scala 971:30]
  wire  tlb_data_register_io_tlb_read_data_v_1; // @[myCPU.scala 971:30]
  wire [18:0] tlb_data_register_io_tlb_write_data_vaddr; // @[myCPU.scala 971:30]
  wire [7:0] tlb_data_register_io_tlb_write_data_asid; // @[myCPU.scala 971:30]
  wire  tlb_data_register_io_tlb_write_data_g; // @[myCPU.scala 971:30]
  wire [19:0] tlb_data_register_io_tlb_write_data_paddr_0; // @[myCPU.scala 971:30]
  wire [19:0] tlb_data_register_io_tlb_write_data_paddr_1; // @[myCPU.scala 971:30]
  wire [2:0] tlb_data_register_io_tlb_write_data_c_0; // @[myCPU.scala 971:30]
  wire [2:0] tlb_data_register_io_tlb_write_data_c_1; // @[myCPU.scala 971:30]
  wire  tlb_data_register_io_tlb_write_data_d_0; // @[myCPU.scala 971:30]
  wire  tlb_data_register_io_tlb_write_data_d_1; // @[myCPU.scala 971:30]
  wire  tlb_data_register_io_tlb_write_data_v_0; // @[myCPU.scala 971:30]
  wire  tlb_data_register_io_tlb_write_data_v_1; // @[myCPU.scala 971:30]
  wire  _T_2 = ~resetn; // @[myCPU.scala 106:41]
  wire  stage_fec_2_inst_jump = inst_sram_rdata_L[33]; // @[myCPU.scala 159:45]
  wire  stage_fec_2_inst_branch = inst_sram_rdata_L[32]; // @[myCPU.scala 160:47]
  reg  pre_decoder_branchD_flag; // @[myCPU.scala 162:44]
  reg [5:0] pre_decoder_branchdata; // @[myCPU.scala 163:43]
  reg  pre_decoder_jump; // @[myCPU.scala 164:40]
  reg  pre_decoder_jr; // @[myCPU.scala 165:40]
  wire  _PCSrcD_T_1 = _cfu_io_StallD; // @[myCPU.scala 179:66]
  wire  _PCSrcD_T_3 = _br_io_exe; // @[myCPU.scala 179:85]
  wire [6:0] PCBranchD_lo = {_if2id_io_InstrD[15],_if2id_io_InstrD[15],_if2id_io_InstrD[15],_if2id_io_InstrD[15],
    _if2id_io_InstrD[15],_if2id_io_InstrD[15],_if2id_io_InstrD[15]}; // @[Cat.scala 31:58]
  wire [31:0] _PCBranchD_T_16 = {_if2id_io_InstrD[15],_if2id_io_InstrD[15],_if2id_io_InstrD[15],_if2id_io_InstrD[15],
    _if2id_io_InstrD[15],_if2id_io_InstrD[15],_if2id_io_InstrD[15],PCBranchD_lo,_if2id_io_InstrD[15:0],2'h0}; // @[Cat.scala 31:58]
  wire [31:0] PCBranchD = _PCBranchD_T_16 + _if2id_io_PCPlus4D; // @[myCPU.scala 180:98]
  wire [31:0] _PCJumpD_T_3 = {_if2id_io_PCPlus4D[31:28],_if2id_io_InstrD[25:0],2'h0}; // @[Cat.scala 31:58]
  reg [31:0] resultE2M_Reg; // @[myCPU.scala 928:32]
  reg [31:0] ResultM2_Reg; // @[myCPU.scala 988:29]
  wire [31:0] _BranchRsD_T_2 = _cfu_io_ForwardAD[1] ? ResultM2_Reg : _regfile_io_RD1; // @[myCPU.scala 739:61]
  wire [31:0] BranchRsD = _cfu_io_ForwardAD[0] ? resultE2M_Reg : _BranchRsD_T_2; // @[myCPU.scala 739:20]
  wire [31:0] PCJumpD = pre_decoder_jr ? BranchRsD : _PCJumpD_T_3; // @[myCPU.scala 181:24]
  wire [4:0] RdD = _if2id_io_InstrD[15:11]; // @[myCPU.scala 184:27]
  wire [16:0] _ImmD_T_3 = {1'h0,_if2id_io_InstrD[15:0]}; // @[Cat.scala 31:58]
  wire [7:0] ImmD_lo = {_if2id_io_InstrD[15],_if2id_io_InstrD[15],_if2id_io_InstrD[15],_if2id_io_InstrD[15],
    _if2id_io_InstrD[15],_if2id_io_InstrD[15],_if2id_io_InstrD[15],_if2id_io_InstrD[15]}; // @[Cat.scala 31:58]
  wire [31:0] _ImmD_T_23 = {_if2id_io_InstrD[15],_if2id_io_InstrD[15],_if2id_io_InstrD[15],_if2id_io_InstrD[15],
    _if2id_io_InstrD[15],_if2id_io_InstrD[15],_if2id_io_InstrD[15],_if2id_io_InstrD[15],ImmD_lo,_if2id_io_InstrD[15:0]}; // @[Cat.scala 31:58]
  wire [2:0] Write_WriteCP0Sel0 = _if2id_io_InstrD[2:0]; // @[myCPU.scala 187:37]
  reg [31:0] PCW_Reg; // @[myCPU.scala 273:26]
  reg  slot_Reg; // @[myCPU.scala 274:27]
  reg [1:0] branchjump_Jr_Reg; // @[myCPU.scala 275:36]
  wire  _PCW_Reg_T = _mem22wb_io_PCW != 32'h0; // @[myCPU.scala 277:36]
  reg [31:0] reg_pc; // @[myCPU.scala 283:25]
  reg  wb_exception; // @[myCPU.scala 602:27]
  wire  RegWriteW = wb_exception ? 1'h0 : _mem22wb_io_RegWriteW_Out; // @[myCPU.scala 1115:21]
  wire [3:0] _debug_wb_rf_wen_T_2 = RegWriteW ? 4'hf : 4'h0; // @[myCPU.scala 286:62]
  reg [31:0] pc_next_wait; // @[myCPU.scala 324:31]
  wire  ready_to_branch = fifo_io_point_write_en; // @[myCPU.scala 326:31 555:21]
  reg  commit_bru_reg; // @[myCPU.scala 380:30]
  reg  stage_fec_2_stall_reg; // @[myCPU.scala 490:40]
  reg  stage_fec_2_valid; // @[myCPU.scala 461:36]
  wire  _stage_fec_2_branch_answer_T_7 = _cp0_io_exception; // @[myCPU.scala 493:209]
  wire  _stage_fec_2_branch_answer_T_8 = ~_cp0_io_exception; // @[myCPU.scala 493:190]
  wire  stage_fec_2_branch_answer = commit_bru_reg & branch_prediction_with_blockram_io_pre_L & (stage_fec_2_inst_branch
     | stage_fec_2_inst_jump) & branch_prediction_with_blockram_io_btb_hit_0 & stage_fec_2_stall_reg & stage_fec_2_valid
     & ~_cp0_io_exception; // @[myCPU.scala 493:187]
  wire  _pc_next_wait_T = ready_to_branch | stage_fec_2_branch_answer; // @[myCPU.scala 327:41]
  wire [31:0] _PC_nextD_T_2 = _PCSrcD_T_3 ? PCBranchD : _if2id_io_PCPlus8D; // @[Mux.scala 101:16]
  wire [31:0] PC_nextD = pre_decoder_jump ? PCJumpD : _PC_nextD_T_2; // @[Mux.scala 101:16]
  wire [31:0] stage_fec_2_pre_target_0 = branch_prediction_with_blockram_io_pre_target_L; // @[myCPU.scala 466:38 482:31]
  wire [31:0] stage_fec_1_pc = stage_fec_1_pc_L_io_out_pc_value_out; // @[myCPU.scala 156:26 431:20]
  wire [31:0] _stage_fec_1_pc_next_T_1 = stage_fec_1_pc + 32'h4; // @[myCPU.scala 398:93]
  wire [31:0] stage_fec_1_pc_next = stage_fec_2_branch_answer ? stage_fec_2_pre_target_0 : _stage_fec_1_pc_next_T_1; // @[myCPU.scala 398:31]
  wire [31:0] Pc_Next_normal = fifo_io_point_write_en ? PC_nextD : stage_fec_1_pc_next; // @[myCPU.scala 731:26]
  reg  pc_req_wait; // @[myCPU.scala 328:30]
  wire  _T_4 = ~inst_sram_en; // @[myCPU.scala 332:10]
  wire  _GEN_0 = pc_req_wait & inst_sram_en | _stage_fec_2_branch_answer_T_7 | ready_to_branch & inst_sram_en ? 1'h0 :
    pc_req_wait; // @[myCPU.scala 334:119 335:21 337:21]
  reg [31:0] exception_Pc_reg; // @[myCPU.scala 341:35]
  reg  returnPc_req_wait; // @[myCPU.scala 344:36]
  wire  _GEN_2 = returnPc_req_wait & inst_sram_en ? 1'h0 : returnPc_req_wait; // @[myCPU.scala 349:54 350:27 352:27]
  wire [31:0] _Pc_Next_T_1 = pc_req_wait ? pc_next_wait : Pc_Next_normal; // @[myCPU.scala 359:140]
  wire [31:0] _Pc_Next_T_2 = ready_to_branch ? Pc_Next_normal : _Pc_Next_T_1; // @[myCPU.scala 359:105]
  wire [31:0] _Pc_Next_T_3 = returnPc_req_wait ? exception_Pc_reg : _Pc_Next_T_2; // @[myCPU.scala 359:66]
  wire [31:0] Pc_Next = _stage_fec_2_branch_answer_T_7 ? _cp0_io_return_pc : _Pc_Next_T_3; // @[myCPU.scala 359:19]
  reg  commit_cache_reg; // @[myCPU.scala 379:32]
  wire  _commit_cache_reg_T = _cfu_io_StallE; // @[myCPU.scala 381:40]
  reg  stage_fec_1_valid; // @[myCPU.scala 440:36]
  wire  _access_stage1_sram_valid_T_1 = fifo_io_empty; // @[myCPU.scala 442:97]
  wire  _access_stage1_sram_valid_T_9 = ready_to_branch & (~fifo_io_empty | fifo_io_empty & inst_write_en != 2'h0) |
    fifo_io_point_flush; // @[myCPU.scala 442:161]
  wire  access_stage1_sram_valid = ~(ready_to_branch & (~fifo_io_empty | fifo_io_empty & inst_write_en != 2'h0) |
    fifo_io_point_flush) & _stage_fec_2_branch_answer_T_8; // @[myCPU.scala 442:196]
  wire  _stage_fec_1_valid_T_1 = ready_to_branch ? access_stage1_sram_valid : stage_fec_1_valid; // @[myCPU.scala 444:55]
  reg [6:0] stage_fec_2_bht_0; // @[myCPU.scala 464:35]
  reg [3:0] stage_fec_2_hascode_0; // @[myCPU.scala 468:39]
  wire  stage_fec_2_hascode_0_num_array_0 = ^branch_prediction_with_blockram_io_pc[7:4]; // @[macros.scala 389:45]
  wire  stage_fec_2_hascode_0_num_array_1 = ^branch_prediction_with_blockram_io_pc[11:8]; // @[macros.scala 389:45]
  wire  stage_fec_2_hascode_0_num_array_2 = ^branch_prediction_with_blockram_io_pc[15:12]; // @[macros.scala 389:45]
  wire  stage_fec_2_hascode_0_num_array_3 = ^branch_prediction_with_blockram_io_pc[19:16]; // @[macros.scala 389:45]
  wire [3:0] _stage_fec_2_hascode_0_T_1 = {stage_fec_2_hascode_0_num_array_3,stage_fec_2_hascode_0_num_array_2,
    stage_fec_2_hascode_0_num_array_1,stage_fec_2_hascode_0_num_array_0}; // @[macros.scala 391:13]
  wire  _stage_fec_2_data_valid_T = ~fifo_io_empty; // @[myCPU.scala 511:88]
  wire [5:0] opD = inst_sram_rdata_L[31:26]; // @[myCPU.scala 108:24]
  wire [5:0] FunctD = inst_sram_rdata_L[5:0]; // @[myCPU.scala 110:27]
  wire  _T_31 = 6'h0 == opD & (6'h9 == FunctD | 6'h8 == FunctD); // @[Mux.scala 81:58]
  wire [6:0] stage_fec_2_lookup_data_0 = branch_prediction_with_blockram_io_lookup_data_0; // @[myCPU.scala 469:40 471:29]
  wire [1:0] stage_fec_2_pht_0 = branch_prediction_with_blockram_io_out_L; // @[myCPU.scala 465:32 478:24]
  wire [108:0] lo = {stage_fec_2_pht_0,stage_fec_2_pre_target_0,stage_fec_2_hascode_0,stage_fec_2_lookup_data_0,
    inst_sram_rdata_L[31:0],stage_fec_2_pc_L_io_out_pc_value_out}; // @[Cat.scala 31:58]
  wire [26:0] hi = {inst_tlb_exception,_T_31,inst_sram_rdata_L[39:32],branch_prediction_with_blockram_io_pht_out,
    stage_fec_2_branch_answer,stage_fec_2_bht_0}; // @[Cat.scala 31:58]
  wire  _T_35 = _cfu_io_StallF; // @[myCPU.scala 535:51]
  wire  _pre_decoder_branchD_flag_T = _cfu_io_FlushD; // @[myCPU.scala 560:52]
  reg  InDelaySlotF; // @[myCPU.scala 566:31]
  wire  _T_54 = pre_decoder_branchD_flag | pre_decoder_jump; // @[myCPU.scala 567:43]
  wire  _GEN_6 = _T_35 ? 1'h0 : InDelaySlotF; // @[myCPU.scala 569:38 570:22 572:22]
  wire  __if2id_io_InstrF_T = _cu_io1_BadInstrD; // @[myCPU.scala 584:52]
  wire  __if2id_io_InstrF_T_1 = _cu_io1_SysCallD; // @[myCPU.scala 584:79]
  wire  __if2id_io_InstrF_T_3 = _cu_io1_BreakD; // @[myCPU.scala 584:102]
  wire  __if2id_io_InstrF_T_5 = _cu_io1_EretD; // @[myCPU.scala 585:23]
  reg  id_exception; // @[myCPU.scala 590:27]
  reg  ex_exception; // @[myCPU.scala 593:27]
  wire  _ex_exception_T = _cfu_io_FlushE; // @[myCPU.scala 594:36]
  reg  mem_exception; // @[myCPU.scala 596:28]
  wire  _mem_exception_T = _cfu_io_FlushM; // @[myCPU.scala 597:37]
  wire  _mem_exception_T_1 = _cfu_io_StallM; // @[myCPU.scala 597:67]
  reg  mem2_exception; // @[myCPU.scala 599:29]
  wire  _mem2_exception_T = _cfu_io_FlushM2; // @[myCPU.scala 600:39]
  wire  _mem2_exception_T_1 = _cfu_io_StallM2; // @[myCPU.scala 600:70]
  wire  _wb_exception_T = _cfu_io_FlushW; // @[myCPU.scala 603:36]
  wire  _wb_exception_T_1 = _cfu_io_StallW; // @[myCPU.scala 603:66]
  reg  id_true_branch_state; // @[myCPU.scala 649:35]
  reg  inst_tlb_exceptionE; // @[myCPU.scala 679:34]
  wire  target_neq_branchD = id_bru_state_io_out_target_pc != PCBranchD; // @[myCPU.scala 693:62]
  wire  target_neq_jumpD = id_bru_state_io_out_target_pc != PCJumpD; // @[myCPU.scala 694:62]
  wire  target_addr_error = pre_decoder_jump & target_neq_jumpD | _PCSrcD_T_3 & target_neq_branchD; // @[myCPU.scala 696:75]
  wire  _T_61 = pre_decoder_jump | _PCSrcD_T_3; // @[myCPU.scala 699:88]
  wire [31:0] _Pc_targetD_T_2 = pre_decoder_jump ? PCJumpD : 32'h0; // @[Mux.scala 101:16]
  reg  true_branch_stateE; // @[myCPU.scala 709:37]
  wire [1:0] _pht_tobeE_T_1 = true_branch_stateE ? 2'h3 : 2'h2; // @[macros.scala 410:30]
  wire [1:0] _pht_tobeE_T_2 = true_branch_stateE ? 2'h2 : 2'h0; // @[macros.scala 411:32]
  wire [1:0] _pht_tobeE_T_3 = true_branch_stateE ? 2'h3 : 2'h1; // @[macros.scala 412:30]
  wire [1:0] _pht_tobeE_T_5 = 2'h3 == ex_bru_state_io_out_pht ? _pht_tobeE_T_1 : {{1'd0}, true_branch_stateE}; // @[Mux.scala 81:58]
  wire [1:0] _pht_tobeE_T_7 = 2'h1 == ex_bru_state_io_out_pht ? _pht_tobeE_T_2 : _pht_tobeE_T_5; // @[Mux.scala 81:58]
  wire [1:0] pht_tobeE = 2'h2 == ex_bru_state_io_out_pht ? _pht_tobeE_T_3 : _pht_tobeE_T_7; // @[Mux.scala 81:58]
  wire [7:0] _pht_lookup_value_tobeE_T_2 = {ex_bru_state_io_out_pht_lookup_value[7:2],pht_tobeE}; // @[Cat.scala 31:58]
  wire [7:0] _pht_lookup_value_tobeE_T_5 = {ex_bru_state_io_out_pht_lookup_value[7:4],pht_tobeE,
    ex_bru_state_io_out_pht_lookup_value[1:0]}; // @[Cat.scala 31:58]
  wire [7:0] _pht_lookup_value_tobeE_T_8 = {ex_bru_state_io_out_pht_lookup_value[7:6],pht_tobeE,
    ex_bru_state_io_out_pht_lookup_value[3:0]}; // @[Cat.scala 31:58]
  wire [7:0] _pht_lookup_value_tobeE_T_10 = {pht_tobeE,ex_bru_state_io_out_pht_lookup_value[5:0]}; // @[Cat.scala 31:58]
  wire [7:0] _pht_lookup_value_tobeE_T_12 = 2'h1 == ex_bru_state_io_out_lookup_data[1:0] ? _pht_lookup_value_tobeE_T_5
     : _pht_lookup_value_tobeE_T_2; // @[Mux.scala 81:58]
  wire [7:0] _pht_lookup_value_tobeE_T_14 = 2'h2 == ex_bru_state_io_out_lookup_data[1:0] ? _pht_lookup_value_tobeE_T_8
     : _pht_lookup_value_tobeE_T_12; // @[Mux.scala 81:58]
  wire [31:0] _BranchRtD_T_2 = _cfu_io_ForwardBD[1] ? ResultM2_Reg : _regfile_io_RD2; // @[myCPU.scala 741:61]
  wire  _ExceptionTypeD_Out_T_1 = _if2id_io_PCD[1:0] != 2'h0; // @[myCPU.scala 743:29]
  wire [20:0] _ExceptionTypeD_Out_T_4 = _ExceptionTypeD_Out_T_1 ? 21'h100000 : 21'h0; // @[Mux.scala 27:73]
  wire [3:0] _ExceptionTypeD_Out_T_5 = _if2id_io_ExceptionTypeD_Out[0] ? 4'h8 : 4'h0; // @[Mux.scala 27:73]
  wire [2:0] _ExceptionTypeD_Out_T_6 = _if2id_io_ExceptionTypeD_Out[1] ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [20:0] _GEN_16 = {{17'd0}, _ExceptionTypeD_Out_T_5}; // @[Mux.scala 27:73]
  wire [20:0] _ExceptionTypeD_Out_T_7 = _ExceptionTypeD_Out_T_4 | _GEN_16; // @[Mux.scala 27:73]
  wire [20:0] _GEN_17 = {{18'd0}, _ExceptionTypeD_Out_T_6}; // @[Mux.scala 27:73]
  wire [20:0] _ExceptionTypeD_Out_T_8 = _ExceptionTypeD_Out_T_7 | _GEN_17; // @[Mux.scala 27:73]
  reg [5:0] int_instanceE; // @[myCPU.scala 751:33]
  reg [5:0] int_instanceM; // @[myCPU.scala 752:33]
  reg [5:0] int_instanceM2; // @[myCPU.scala 753:33]
  reg [5:0] int_instanceW; // @[myCPU.scala 754:33]
  wire  _int_with_timer_int_T_1 = _cp0_io_timer_int_has | ext_int[5]; // @[myCPU.scala 756:56]
  wire [5:0] int_with_timer_int = {_int_with_timer_int_T_1,ext_int[4:0]}; // @[Cat.scala 31:58]
  wire [5:0] __id2ex_io_ExceptionTypeD_T = int_with_timer_int & _cp0_io_cp0_status; // @[myCPU.scala 767:59]
  wire [31:0] ExceptionTypeD_Out = {{11'd0}, _ExceptionTypeD_Out_T_8}; // @[myCPU.scala 171:34 742:24]
  wire [10:0] __id2ex_io_ExceptionTypeD_T_6 = __if2id_io_InstrF_T ? 11'h400 : 11'h0; // @[myCPU.scala 768:13]
  wire [8:0] __id2ex_io_ExceptionTypeD_T_8 = __if2id_io_InstrF_T_1 ? 9'h100 : 9'h0; // @[myCPU.scala 769:13]
  wire [10:0] _GEN_18 = {{2'd0}, __id2ex_io_ExceptionTypeD_T_8}; // @[myCPU.scala 768:59]
  wire [10:0] __id2ex_io_ExceptionTypeD_T_9 = __id2ex_io_ExceptionTypeD_T_6 | _GEN_18; // @[myCPU.scala 768:59]
  wire [9:0] __id2ex_io_ExceptionTypeD_T_11 = __if2id_io_InstrF_T_3 ? 10'h200 : 10'h0; // @[myCPU.scala 770:13]
  wire [10:0] _GEN_19 = {{1'd0}, __id2ex_io_ExceptionTypeD_T_11}; // @[myCPU.scala 769:59]
  wire [10:0] __id2ex_io_ExceptionTypeD_T_12 = __id2ex_io_ExceptionTypeD_T_9 | _GEN_19; // @[myCPU.scala 769:59]
  wire [31:0] __id2ex_io_ExceptionTypeD_T_14 = __if2id_io_InstrF_T_5 ? 32'h80000000 : 32'h0; // @[myCPU.scala 771:13]
  wire [31:0] _GEN_20 = {{21'd0}, __id2ex_io_ExceptionTypeD_T_12}; // @[myCPU.scala 770:59]
  wire [31:0] __id2ex_io_ExceptionTypeD_T_15 = _GEN_20 | __id2ex_io_ExceptionTypeD_T_14; // @[myCPU.scala 770:59]
  wire [31:0] __id2ex_io_ExceptionTypeD_T_16 = ExceptionTypeD_Out == 32'h0 ? __id2ex_io_ExceptionTypeD_T_15 :
    ExceptionTypeD_Out; // @[myCPU.scala 767:135]
  wire [4:0] __id2ex_io_ReadCP0AddrD_T_5 = _cu_io1_Tlb_Control[0] ? 5'h0 : RdD; // @[Mux.scala 101:16]
  wire [4:0] __id2ex_io_ReadCP0AddrD_T_6 = _cu_io1_Tlb_Control[1] ? 5'h0 : __id2ex_io_ReadCP0AddrD_T_5; // @[Mux.scala 101:16]
  wire [4:0] __id2ex_io_ReadCP0AddrD_T_7 = _cu_io1_Tlb_Control[2] ? 5'ha : __id2ex_io_ReadCP0AddrD_T_6; // @[Mux.scala 101:16]
  reg  inst_tlb_exceptionM; // @[myCPU.scala 806:34]
  wire [31:0] ResultW = _mem22wb_io_ResultW; // @[myCPU.scala 1114:15 270:26]
  wire [31:0] _RD1ForWardE_p_T_1 = 2'h1 == _cfu_io_ForwardAE ? ResultW : _id2ex_io_RD1E; // @[Mux.scala 81:58]
  wire [31:0] _RD1ForWardE_p_T_3 = 2'h2 == _cfu_io_ForwardAE ? resultE2M_Reg : _RD1ForWardE_p_T_1; // @[Mux.scala 81:58]
  wire [31:0] RD1ForWardE_p = 2'h3 == _cfu_io_ForwardAE ? ResultM2_Reg : _RD1ForWardE_p_T_3; // @[Mux.scala 81:58]
  wire [31:0] _RD2ForWardE_p_T_1 = 2'h1 == _cfu_io_ForwardBE ? ResultW : _id2ex_io_RD2E; // @[Mux.scala 81:58]
  wire [31:0] _RD2ForWardE_p_T_3 = 2'h2 == _cfu_io_ForwardBE ? resultE2M_Reg : _RD2ForWardE_p_T_1; // @[Mux.scala 81:58]
  wire [31:0] RD2ForWardE_p = 2'h3 == _cfu_io_ForwardBE ? ResultM2_Reg : _RD2ForWardE_p_T_3; // @[Mux.scala 81:58]
  reg [31:0] RD1ForWardE_r; // @[myCPU.scala 811:34]
  reg [31:0] RD2ForWardE_r; // @[myCPU.scala 812:34]
  reg  Forward_Lock1E; // @[myCPU.scala 813:34]
  reg  Forward_Lock2E; // @[myCPU.scala 814:34]
  wire [31:0] _Forward_CP0_data_T_1 = 2'h1 == _cfu_io_ForwardCP0E ? _ex2mem_io_WriteCP0HiLoDataM : _cp0_io_cp0_read_data
    ; // @[Mux.scala 81:58]
  wire [31:0] Forward_CP0_data = 2'h2 == _cfu_io_ForwardCP0E ? _mem2mem2_io_WriteCP0HiLoDataM : _Forward_CP0_data_T_1; // @[Mux.scala 81:58]
  wire [31:0] RD1ForWardE = Forward_Lock1E ? RD1ForWardE_r : RD1ForWardE_p; // @[myCPU.scala 819:23]
  wire [31:0] RD2ForWardE = Forward_Lock2E ? RD2ForWardE_r : RD2ForWardE_p; // @[myCPU.scala 820:23]
  wire  _Forward_Lock1E_T = _ex2mem_io_MemToRegM; // @[myCPU.scala 826:54]
  wire  _Forward_Lock1E_T_1 = _mem2mem2_io_MemToRegM; // @[myCPU.scala 826:87]
  wire  _Forward_Lock1E_T_3 = ~(_ex2mem_io_MemToRegM | _mem2mem2_io_MemToRegM); // @[myCPU.scala 826:31]
  wire [31:0] Inst_badvaddrE = _id2ex_io_ExceptionTypeE_Out[31] ? Forward_CP0_data : _id2ex_io_BadVaddrE; // @[myCPU.scala 836:29]
  wire [4:0] _WriteRegE_T_1 = 2'h1 == _id2ex_io2_RegDstE ? _id2ex_io_RdE : _id2ex_io_RtE; // @[Mux.scala 81:58]
  wire [4:0] _WriteRegE_T_3 = 2'h2 == _id2ex_io2_RegDstE ? 5'h1f : _WriteRegE_T_1; // @[Mux.scala 81:58]
  wire  _WriteCP0HiLoDataE_T_1 = _id2ex_io2_CP0WriteE; // @[myCPU.scala 841:30]
  wire [31:0] _WriteCP0HiLoDataE_T_2 = _WriteCP0HiLoDataE_T_1 ? RD2ForWardE : 32'h0; // @[myCPU.scala 840:79]
  wire [31:0] WriteCP0HiLoDataE = _id2ex_io2_HiLoWriteE != 2'h0 ? RD1ForWardE : _WriteCP0HiLoDataE_T_2; // @[myCPU.scala 840:32]
  wire [31:0] _Src1E_T_3 = {27'h0,_id2ex_io_ImmE[10:6]}; // @[Cat.scala 31:58]
  wire  CP0ToRegE = _id2ex_io_ExceptionTypeE_Out == 32'h0 & _id2ex_io_CP0ToRegE_Out; // @[myCPU.scala 844:24]
  wire [2:0] _muldiv_io_ctrl_hi = {_id2ex_io2_ALUCtrlE[21],_id2ex_io2_ALUCtrlE[9:8]}; // @[Cat.scala 31:58]
  wire  __dmemreq_io_en_T_3 = _addr_cal_io_d_unaligned; // @[myCPU.scala 863:71]
  wire  __dmemreq_io_en_T_6 = ~_addr_cal_io_d_unaligned & _commit_cache_reg_T; // @[myCPU.scala 863:78]
  wire [31:0] __ex2mem_io_HiLoOutE_T_2 = 2'h1 == _cfu_io_ForwardHE ? _mem22wb_io_LoInW : _hilo_io_lo_o; // @[Mux.scala 81:58]
  wire [31:0] __ex2mem_io_HiLoOutE_T_4 = 2'h2 == _cfu_io_ForwardHE ? _ex2mem_io_LoInM : __ex2mem_io_HiLoOutE_T_2; // @[Mux.scala 81:58]
  wire [31:0] __ex2mem_io_HiLoOutE_T_6 = 2'h3 == _cfu_io_ForwardHE ? _mem2mem2_io_LoInM : __ex2mem_io_HiLoOutE_T_4; // @[Mux.scala 81:58]
  wire [31:0] __ex2mem_io_HiLoOutE_T_9 = 2'h1 == _cfu_io_ForwardHE ? _mem22wb_io_HiInW : _hilo_io_hi_o; // @[Mux.scala 81:58]
  wire [31:0] __ex2mem_io_HiLoOutE_T_11 = 2'h2 == _cfu_io_ForwardHE ? _ex2mem_io_HiInM : __ex2mem_io_HiLoOutE_T_9; // @[Mux.scala 81:58]
  wire [31:0] __ex2mem_io_HiLoOutE_T_13 = 2'h3 == _cfu_io_ForwardHE ? _mem2mem2_io_HiInM : __ex2mem_io_HiLoOutE_T_11; // @[Mux.scala 81:58]
  wire [31:0] __ex2mem_io_HiLoOutE_T_14 = _id2ex_io2_HiLoToRegE[0] ? __ex2mem_io_HiLoOutE_T_6 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] __ex2mem_io_HiLoOutE_T_15 = _id2ex_io2_HiLoToRegE[1] ? __ex2mem_io_HiLoOutE_T_13 : 32'h0; // @[Mux.scala 27:73]
  wire  _temp_exceptionE_T_2 = _id2ex_io2_MemToRegE; // @[myCPU.scala 882:70]
  wire [4:0] _temp_exceptionE_T_4 = __dmemreq_io_en_T_3 & _id2ex_io2_MemToRegE ? 5'h10 : 5'h0; // @[myCPU.scala 882:13]
  wire  _temp_exceptionE_T_6 = _id2ex_io2_MemWriteE; // @[myCPU.scala 883:70]
  wire [5:0] _temp_exceptionE_T_8 = __dmemreq_io_en_T_3 & _id2ex_io2_MemWriteE ? 6'h20 : 6'h0; // @[myCPU.scala 883:13]
  wire [5:0] _GEN_21 = {{1'd0}, _temp_exceptionE_T_4}; // @[myCPU.scala 882:101]
  wire [5:0] _temp_exceptionE_T_9 = _GEN_21 | _temp_exceptionE_T_8; // @[myCPU.scala 882:101]
  wire [12:0] _temp_exceptionE_T_11 = _alu_io_overflow ? 13'h1000 : 13'h0; // @[myCPU.scala 884:13]
  wire [12:0] _GEN_22 = {{7'd0}, _temp_exceptionE_T_9}; // @[myCPU.scala 883:101]
  wire [12:0] _temp_exceptionE_T_12 = _GEN_22 | _temp_exceptionE_T_11; // @[myCPU.scala 883:101]
  wire [31:0] temp_exceptionE = _id2ex_io_ExceptionTypeE_Out != 32'h0 ? _id2ex_io_ExceptionTypeE_Out : {{19'd0},
    _temp_exceptionE_T_12}; // @[myCPU.scala 881:30]
  wire  _Forward_for_epc_T = _ex2mem_io_CP0WriteM; // @[myCPU.scala 889:52]
  wire  _Forward_for_epc_T_5 = _mem2mem2_io_CP0WriteM & _mem2mem2_io_WriteCP0AddrM == 5'he; // @[myCPU.scala 890:39]
  wire [31:0] _Forward_for_epc_T_6 = _Forward_for_epc_T_5 ? _mem2mem2_io_WriteCP0HiLoDataM : _cp0_io_epc; // @[myCPU.scala 889:134]
  wire [31:0] Forward_for_epc = _ex2mem_io_CP0WriteM & _ex2mem_io_WriteCP0AddrM == 5'he ? _ex2mem_io_WriteCP0HiLoDataM
     : _Forward_for_epc_T_6; // @[myCPU.scala 889:30]
  wire  _BadVAddrE_T_8 = _id2ex_io_ExceptionTypeE_Out[31] & Forward_for_epc[1:0] != 2'h0; // @[myCPU.scala 892:175]
  wire [31:0] _BadVAddrE_T_9 = _id2ex_io_ExceptionTypeE_Out[31] & Forward_for_epc[1:0] != 2'h0 ? Forward_for_epc :
    Inst_badvaddrE; // @[myCPU.scala 892:141]
  wire [20:0] __ex2mem_io_ExceptionTypeE_T_4 = _BadVAddrE_T_8 ? 21'h100000 : 21'h0; // @[myCPU.scala 896:39]
  wire [31:0] _GEN_23 = {{11'd0}, __ex2mem_io_ExceptionTypeE_T_4}; // @[myCPU.scala 896:127]
  wire  _resultE_T_1 = _id2ex_io2_HiLoToRegE != 2'h0; // @[myCPU.scala 923:32]
  wire  _resultE_T_2 = _id2ex_io2_LinkE; // @[myCPU.scala 924:25]
  wire [31:0] _resultE_T_4 = _id2ex_io2_ALUCtrlE[21] ? _muldiv_io_lo : _alu_io_result; // @[Mux.scala 101:16]
  wire [31:0] _resultE_T_5 = _resultE_T_2 ? _id2ex_io2_PCPlus8E : _resultE_T_4; // @[Mux.scala 101:16]
  wire  _tlb_searched_index_value_T = ~tlb_search_hit; // @[myCPU.scala 986:33]
  wire [31:0] tlb_searched_index_value = {_tlb_searched_index_value_T,27'h0,tlb_search_index}; // @[Cat.scala 31:58]
  wire [6:0] _ExceptionM_T_2 = _Forward_Lock1E_T ? 7'h8 : 7'h40; // @[myCPU.scala 993:33]
  wire [7:0] _ExceptionM_T_5 = _Forward_Lock1E_T ? 8'h4 : 8'h80; // @[myCPU.scala 994:33]
  wire [6:0] _ExceptionM_T_7 = data_tlb_exception[0] ? _ExceptionM_T_2 : 7'h0; // @[Mux.scala 27:73]
  wire [7:0] _ExceptionM_T_8 = data_tlb_exception[1] ? _ExceptionM_T_5 : 8'h0; // @[Mux.scala 27:73]
  wire [1:0] _ExceptionM_T_9 = data_tlb_exception[2] ? 2'h2 : 2'h0; // @[Mux.scala 27:73]
  wire [7:0] _GEN_24 = {{1'd0}, _ExceptionM_T_7}; // @[Mux.scala 27:73]
  wire [7:0] _ExceptionM_T_10 = _GEN_24 | _ExceptionM_T_8; // @[Mux.scala 27:73]
  wire [7:0] _GEN_25 = {{6'd0}, _ExceptionM_T_9}; // @[Mux.scala 27:73]
  wire [7:0] _ExceptionM_T_11 = _ExceptionM_T_10 | _GEN_25; // @[Mux.scala 27:73]
  wire  __mem2mem2_io_CP0WriteE_T_2 = _Forward_for_epc_T | _ex2mem_io_Tlb_ControlM[2]; // @[myCPU.scala 1002:55]
  wire  __mem2mem2_io_WriteCP0HiLoDataE_T = data_tlb_exception != 3'h0; // @[myCPU.scala 1005:25]
  wire [31:0] __mem2mem2_io_WriteCP0HiLoDataE_T_2 = {_ex2mem_io_PhyAddrM[31:13],5'h0,_cp0_io_asid}; // @[Cat.scala 31:58]
  wire [31:0] __mem2mem2_io_WriteCP0HiLoDataE_T_5 = {_ex2mem_io_PCM[31:13],5'h0,_cp0_io_asid}; // @[Cat.scala 31:58]
  wire [31:0] __mem2mem2_io_WriteCP0HiLoDataE_T_6 = inst_tlb_exceptionM ? __mem2mem2_io_WriteCP0HiLoDataE_T_5 :
    _ex2mem_io_WriteCP0HiLoDataM; // @[Mux.scala 101:16]
  wire [31:0] __mem2mem2_io_WriteCP0HiLoDataE_T_7 = _ex2mem_io_Tlb_ControlM[2] ? tlb_searched_index_value :
    __mem2mem2_io_WriteCP0HiLoDataE_T_6; // @[Mux.scala 101:16]
  wire  __mem2mem2_io1_WriteCP0AddrE_T_1 = __mem2mem2_io_WriteCP0HiLoDataE_T | inst_tlb_exceptionM; // @[myCPU.scala 1024:64]
  reg  tlb_exception_cp0_writeM2; // @[myCPU.scala 1041:40]
  reg  tlb_exception_co0_writeW; // @[myCPU.scala 1042:40]
  wire [31:0] __mem2mem2_io_BadVAddrE_T_1 = {{20'd0}, _ex2mem_io_ExceptionTypeM_Out[31:20]}; // @[myCPU.scala 1049:117]
  wire  __mem2mem2_io_BadVAddrE_T_4 = ~_ex2mem_io_BadVAddrM[31]; // @[myCPU.scala 1049:160]
  wire  __mem2mem2_io_BadVAddrE_T_7 = __mem2mem2_io_BadVAddrE_T_4 | _ex2mem_io_BadVAddrM[31:30] == 2'h3; // @[myCPU.scala 1050:5]
  wire [31:0] __mem2mem2_io_BadVAddrE_T_9 = __mem2mem2_io_BadVAddrE_T_1[0] & __mem2mem2_io_BadVAddrE_T_7 ?
    _ex2mem_io_PCM : _ex2mem_io_BadVAddrM; // @[myCPU.scala 1049:87]
  wire [31:0] _Mem_withRL_Data_T_25 = {_mem2mem2_io_RtM[31:8],_dmem_io_RD[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _Mem_withRL_Data_T_22 = {_mem2mem2_io_RtM[31:16],_dmem_io_RD[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _Mem_withRL_Data_T_19 = {_mem2mem2_io_RtM[31:24],_dmem_io_RD[31:8]}; // @[Cat.scala 31:58]
  wire [31:0] _Mem_withRL_Data_T_27 = 2'h1 == _mem2mem2_io_PhyAddrM[1:0] ? _Mem_withRL_Data_T_19 : _dmem_io_RD; // @[Mux.scala 81:58]
  wire [31:0] _Mem_withRL_Data_T_29 = 2'h2 == _mem2mem2_io_PhyAddrM[1:0] ? _Mem_withRL_Data_T_22 : _Mem_withRL_Data_T_27
    ; // @[Mux.scala 81:58]
  wire [31:0] _Mem_withRL_Data_T_31 = 2'h3 == _mem2mem2_io_PhyAddrM[1:0] ? _Mem_withRL_Data_T_25 : _Mem_withRL_Data_T_29
    ; // @[Mux.scala 81:58]
  wire [31:0] _Mem_withRL_Data_T_9 = {_dmem_io_RD[23:0],_mem2mem2_io_RtM[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _Mem_withRL_Data_T_6 = {_dmem_io_RD[15:0],_mem2mem2_io_RtM[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _Mem_withRL_Data_T_3 = {_dmem_io_RD[7:0],_mem2mem2_io_RtM[23:0]}; // @[Cat.scala 31:58]
  wire [31:0] _Mem_withRL_Data_T_11 = 2'h0 == _mem2mem2_io_PhyAddrM[1:0] ? _Mem_withRL_Data_T_3 : _dmem_io_RD; // @[Mux.scala 81:58]
  wire [31:0] _Mem_withRL_Data_T_13 = 2'h1 == _mem2mem2_io_PhyAddrM[1:0] ? _Mem_withRL_Data_T_6 : _Mem_withRL_Data_T_11; // @[Mux.scala 81:58]
  wire [31:0] _Mem_withRL_Data_T_15 = 2'h2 == _mem2mem2_io_PhyAddrM[1:0] ? _Mem_withRL_Data_T_9 : _Mem_withRL_Data_T_13; // @[Mux.scala 81:58]
  wire [31:0] _Mem_withRL_Data_T_33 = 2'h2 == _mem2mem2_io_MemRLM ? _Mem_withRL_Data_T_15 : _dmem_io_RD; // @[Mux.scala 81:58]
  wire [31:0] Mem_withRL_Data = 2'h1 == _mem2mem2_io_MemRLM ? _Mem_withRL_Data_T_31 : _Mem_withRL_Data_T_33; // @[Mux.scala 81:58]
  wire  CP0WriteW = wb_exception ? 1'h0 : _mem22wb_io_CP0WriteW; // @[myCPU.scala 1117:25]
  alu _alu ( // @[myCPU.scala 120:22]
    .io_ctrl(_alu_io_ctrl),
    .io_in1(_alu_io_in1),
    .io_in2(_alu_io_in2),
    .io_result(_alu_io_result),
    .io_overflow(_alu_io_overflow)
  );
  br _br ( // @[myCPU.scala 121:22]
    .reset(_br_reset),
    .io_rs(_br_io_rs),
    .io_rt(_br_io_rt),
    .io_branch(_br_io_branch),
    .io_exe(_br_io_exe)
  );
  cfu _cfu ( // @[myCPU.scala 122:22]
    .reset(_cfu_reset),
    .io_Inst_Fifo_Empty(_cfu_io_Inst_Fifo_Empty),
    .io_dmem_calD(_cfu_io_dmem_calD),
    .io_BranchD_Flag(_cfu_io_BranchD_Flag),
    .io_JRD(_cfu_io_JRD),
    .io_CanBranchD(_cfu_io_CanBranchD),
    .io_DivPendingE(_cfu_io_DivPendingE),
    .io_DataPendingM(_cfu_io_DataPendingM),
    .io_InException(_cfu_io_InException),
    .io_WriteRegE(_cfu_io_WriteRegE),
    .io_RegWriteE(_cfu_io_RegWriteE),
    .io_HiLoToRegE(_cfu_io_HiLoToRegE),
    .io_CP0ToRegE(_cfu_io_CP0ToRegE),
    .io_WriteRegM(_cfu_io_WriteRegM),
    .io_MemToRegM(_cfu_io_MemToRegM),
    .io_RegWriteM(_cfu_io_RegWriteM),
    .io_HiLoWriteM(_cfu_io_HiLoWriteM),
    .io_CP0WriteM(_cfu_io_CP0WriteM),
    .io_WriteRegM2(_cfu_io_WriteRegM2),
    .io_MemToRegM2(_cfu_io_MemToRegM2),
    .io_RegWriteM2(_cfu_io_RegWriteM2),
    .io_HiLoWriteM2(_cfu_io_HiLoWriteM2),
    .io_CP0WriteM2(_cfu_io_CP0WriteM2),
    .io_WriteRegW(_cfu_io_WriteRegW),
    .io_RegWriteW(_cfu_io_RegWriteW),
    .io_HiLoWriteW(_cfu_io_HiLoWriteW),
    .io_CP0WriteW(_cfu_io_CP0WriteW),
    .io_ReadCP0AddrE(_cfu_io_ReadCP0AddrE),
    .io_ReadCP0SelE(_cfu_io_ReadCP0SelE),
    .io_WriteCP0AddrM(_cfu_io_WriteCP0AddrM),
    .io_WriteCP0SelM(_cfu_io_WriteCP0SelM),
    .io_WriteCP0AddrM2(_cfu_io_WriteCP0AddrM2),
    .io_WriteCP0SelM2(_cfu_io_WriteCP0SelM2),
    .io_RsD(_cfu_io_RsD),
    .io_RtD(_cfu_io_RtD),
    .io_RsE(_cfu_io_RsE),
    .io_RtE(_cfu_io_RtE),
    .io_StallF(_cfu_io_StallF),
    .io_StallD(_cfu_io_StallD),
    .io_StallE(_cfu_io_StallE),
    .io_StallM(_cfu_io_StallM),
    .io_StallM2(_cfu_io_StallM2),
    .io_StallW(_cfu_io_StallW),
    .io_FlushD(_cfu_io_FlushD),
    .io_FlushE(_cfu_io_FlushE),
    .io_FlushM(_cfu_io_FlushM),
    .io_FlushM2(_cfu_io_FlushM2),
    .io_FlushW(_cfu_io_FlushW),
    .io_ForwardAE(_cfu_io_ForwardAE),
    .io_ForwardBE(_cfu_io_ForwardBE),
    .io_ForwardAD(_cfu_io_ForwardAD),
    .io_ForwardBD(_cfu_io_ForwardBD),
    .io_ForwardHE(_cfu_io_ForwardHE),
    .io_ForwardCP0E(_cfu_io_ForwardCP0E)
  );
  cp0 _cp0 ( // @[myCPU.scala 123:22]
    .clock(_cp0_clock),
    .reset(_cp0_reset),
    .io_cp0_read_addr(_cp0_io_cp0_read_addr),
    .io_cp0_read_sel(_cp0_io_cp0_read_sel),
    .io_cp0_write_addr(_cp0_io_cp0_write_addr),
    .io_cp0_write_sel(_cp0_io_cp0_write_sel),
    .io_cp0_write_data(_cp0_io_cp0_write_data),
    .io_cp0_write_en(_cp0_io_cp0_write_en),
    .io_int_i(_cp0_io_int_i),
    .io_timer_int_has(_cp0_io_timer_int_has),
    .io_pc(_cp0_io_pc),
    .io_mem_bad_vaddr(_cp0_io_mem_bad_vaddr),
    .io_exception_type_i(_cp0_io_exception_type_i),
    .io_in_delayslot(_cp0_io_in_delayslot),
    .io_in_branchjump_jr(_cp0_io_in_branchjump_jr),
    .io_return_pc(_cp0_io_return_pc),
    .io_exception(_cp0_io_exception),
    .io_cp0_read_data(_cp0_io_cp0_read_data),
    .io_epc(_cp0_io_epc),
    .io_cp0_status(_cp0_io_cp0_status),
    .io_Int_able(_cp0_io_Int_able),
    .io_asid(_cp0_io_asid),
    .io_cp0_tlb_read_data_vaddr(_cp0_io_cp0_tlb_read_data_vaddr),
    .io_cp0_tlb_read_data_asid(_cp0_io_cp0_tlb_read_data_asid),
    .io_cp0_tlb_read_data_g(_cp0_io_cp0_tlb_read_data_g),
    .io_cp0_tlb_read_data_paddr_0(_cp0_io_cp0_tlb_read_data_paddr_0),
    .io_cp0_tlb_read_data_paddr_1(_cp0_io_cp0_tlb_read_data_paddr_1),
    .io_cp0_tlb_read_data_c_0(_cp0_io_cp0_tlb_read_data_c_0),
    .io_cp0_tlb_read_data_c_1(_cp0_io_cp0_tlb_read_data_c_1),
    .io_cp0_tlb_read_data_d_0(_cp0_io_cp0_tlb_read_data_d_0),
    .io_cp0_tlb_read_data_d_1(_cp0_io_cp0_tlb_read_data_d_1),
    .io_cp0_tlb_read_data_v_0(_cp0_io_cp0_tlb_read_data_v_0),
    .io_cp0_tlb_read_data_v_1(_cp0_io_cp0_tlb_read_data_v_1),
    .io_cp0_tlb_write_data_vaddr(_cp0_io_cp0_tlb_write_data_vaddr),
    .io_cp0_tlb_write_data_asid(_cp0_io_cp0_tlb_write_data_asid),
    .io_cp0_tlb_write_data_g(_cp0_io_cp0_tlb_write_data_g),
    .io_cp0_tlb_write_data_paddr_0(_cp0_io_cp0_tlb_write_data_paddr_0),
    .io_cp0_tlb_write_data_paddr_1(_cp0_io_cp0_tlb_write_data_paddr_1),
    .io_cp0_tlb_write_data_c_0(_cp0_io_cp0_tlb_write_data_c_0),
    .io_cp0_tlb_write_data_c_1(_cp0_io_cp0_tlb_write_data_c_1),
    .io_cp0_tlb_write_data_d_0(_cp0_io_cp0_tlb_write_data_d_0),
    .io_cp0_tlb_write_data_d_1(_cp0_io_cp0_tlb_write_data_d_1),
    .io_cp0_tlb_write_data_v_0(_cp0_io_cp0_tlb_write_data_v_0),
    .io_cp0_tlb_write_data_v_1(_cp0_io_cp0_tlb_write_data_v_1),
    .io_cp0_tlb_write_en(_cp0_io_cp0_tlb_write_en),
    .io_cp0_index_tlb_write_able(_cp0_io_cp0_index_tlb_write_able)
  );
  cu _cu ( // @[myCPU.scala 124:22]
    .reset(_cu_reset),
    .io1_InstrD(_cu_io1_InstrD),
    .io1_BadInstrD(_cu_io1_BadInstrD),
    .io1_BreakD(_cu_io1_BreakD),
    .io1_SysCallD(_cu_io1_SysCallD),
    .io1_EretD(_cu_io1_EretD),
    .io1_Tlb_Control(_cu_io1_Tlb_Control),
    .io1_commit_cache_ins(_cu_io1_commit_cache_ins),
    .io1_dmem_addr_cal(_cu_io1_dmem_addr_cal),
    .io_RegWriteD(_cu_io_RegWriteD),
    .io_MemToRegD(_cu_io_MemToRegD),
    .io_MemWriteD(_cu_io_MemWriteD),
    .io_ALUCtrlD(_cu_io_ALUCtrlD),
    .io_ALUSrcD(_cu_io_ALUSrcD),
    .io_RegDstD(_cu_io_RegDstD),
    .io_ImmUnsigned(_cu_io_ImmUnsigned),
    .io_LinkD(_cu_io_LinkD),
    .io_HiLoWriteD(_cu_io_HiLoWriteD),
    .io_HiLoToRegD(_cu_io_HiLoToRegD),
    .io_CP0WriteD(_cu_io_CP0WriteD),
    .io_CP0ToRegD(_cu_io_CP0ToRegD),
    .io_LoadUnsignedD(_cu_io_LoadUnsignedD),
    .io_MemWidthD(_cu_io_MemWidthD),
    .io_MemRLD(_cu_io_MemRLD)
  );
  dmem _dmem ( // @[myCPU.scala 125:23]
    .io_data_ok(_dmem_io_data_ok),
    .io_rdata(_dmem_io_rdata),
    .io_Physisc_Address(_dmem_io_Physisc_Address),
    .io_WIDTH(_dmem_io_WIDTH),
    .io_SIGN(_dmem_io_SIGN),
    .io_RD(_dmem_io_RD),
    .io_data_pending(_dmem_io_data_pending)
  );
  dmemreq _dmemreq ( // @[myCPU.scala 126:26]
    .io_en(_dmemreq_io_en),
    .io_MemWriteE(_dmemreq_io_MemWriteE),
    .io_MemToRegE(_dmemreq_io_MemToRegE),
    .io_MemWidthE(_dmemreq_io_MemWidthE),
    .io_VAddrE(_dmemreq_io_VAddrE),
    .io_WriteDataE(_dmemreq_io_WriteDataE),
    .io_memrl(_dmemreq_io_memrl),
    .io_req(_dmemreq_io_req),
    .io_wr(_dmemreq_io_wr),
    .io_size(_dmemreq_io_size),
    .io_addr(_dmemreq_io_addr),
    .io_wdata(_dmemreq_io_wdata),
    .io_wstrb(_dmemreq_io_wstrb)
  );
  ex2mem _ex2mem ( // @[myCPU.scala 127:26]
    .clock(_ex2mem_clock),
    .reset(_ex2mem_reset),
    .io1_RegWriteE(_ex2mem_io1_RegWriteE),
    .io1_MemToRegE(_ex2mem_io1_MemToRegE),
    .io1_LoadUnsignedE(_ex2mem_io1_LoadUnsignedE),
    .io1_MemWidthE(_ex2mem_io1_MemWidthE),
    .io1_HiLoWriteE(_ex2mem_io1_HiLoWriteE),
    .io1_CP0WriteE(_ex2mem_io1_CP0WriteE),
    .io1_WriteCP0AddrE(_ex2mem_io1_WriteCP0AddrE),
    .io1_WriteCP0SelE(_ex2mem_io1_WriteCP0SelE),
    .io1_PCE(_ex2mem_io1_PCE),
    .io1_InDelaySlotE(_ex2mem_io1_InDelaySlotE),
    .io1_MemRLE(_ex2mem_io1_MemRLE),
    .io1_BranchJump_JrE(_ex2mem_io1_BranchJump_JrE),
    .io1_Tlb_Control(_ex2mem_io1_Tlb_Control),
    .io_en(_ex2mem_io_en),
    .io_clr(_ex2mem_io_clr),
    .io_WriteRegE(_ex2mem_io_WriteRegE),
    .io_PhyAddrE(_ex2mem_io_PhyAddrE),
    .io_HiLoOutE(_ex2mem_io_HiLoOutE),
    .io_HiInE(_ex2mem_io_HiInE),
    .io_LoInE(_ex2mem_io_LoInE),
    .io_WriteCP0HiLoDataE(_ex2mem_io_WriteCP0HiLoDataE),
    .io_BadVAddrE(_ex2mem_io_BadVAddrE),
    .io_ExceptionTypeE(_ex2mem_io_ExceptionTypeE),
    .io_RtE(_ex2mem_io_RtE),
    .io_RegWriteM(_ex2mem_io_RegWriteM),
    .io_MemToRegM(_ex2mem_io_MemToRegM),
    .io_WriteRegM(_ex2mem_io_WriteRegM),
    .io_LoadUnsignedM(_ex2mem_io_LoadUnsignedM),
    .io_MemWidthM(_ex2mem_io_MemWidthM),
    .io_PhyAddrM(_ex2mem_io_PhyAddrM),
    .io_HiLoWriteM(_ex2mem_io_HiLoWriteM),
    .io_HiLoOutM(_ex2mem_io_HiLoOutM),
    .io_HiInM(_ex2mem_io_HiInM),
    .io_LoInM(_ex2mem_io_LoInM),
    .io_CP0WriteM(_ex2mem_io_CP0WriteM),
    .io_WriteCP0AddrM(_ex2mem_io_WriteCP0AddrM),
    .io_WriteCP0SelM(_ex2mem_io_WriteCP0SelM),
    .io_WriteCP0HiLoDataM(_ex2mem_io_WriteCP0HiLoDataM),
    .io_PCM(_ex2mem_io_PCM),
    .io_InDelaySlotM(_ex2mem_io_InDelaySlotM),
    .io_BadVAddrM(_ex2mem_io_BadVAddrM),
    .io_ExceptionTypeM_Out(_ex2mem_io_ExceptionTypeM_Out),
    .io_MemRLM(_ex2mem_io_MemRLM),
    .io_RtM(_ex2mem_io_RtM),
    .io_BranchJump_JrM(_ex2mem_io_BranchJump_JrM),
    .io_Tlb_ControlM(_ex2mem_io_Tlb_ControlM)
  );
  ex2mem _mem2mem2 ( // @[myCPU.scala 128:28]
    .clock(_mem2mem2_clock),
    .reset(_mem2mem2_reset),
    .io1_RegWriteE(_mem2mem2_io1_RegWriteE),
    .io1_MemToRegE(_mem2mem2_io1_MemToRegE),
    .io1_LoadUnsignedE(_mem2mem2_io1_LoadUnsignedE),
    .io1_MemWidthE(_mem2mem2_io1_MemWidthE),
    .io1_HiLoWriteE(_mem2mem2_io1_HiLoWriteE),
    .io1_CP0WriteE(_mem2mem2_io1_CP0WriteE),
    .io1_WriteCP0AddrE(_mem2mem2_io1_WriteCP0AddrE),
    .io1_WriteCP0SelE(_mem2mem2_io1_WriteCP0SelE),
    .io1_PCE(_mem2mem2_io1_PCE),
    .io1_InDelaySlotE(_mem2mem2_io1_InDelaySlotE),
    .io1_MemRLE(_mem2mem2_io1_MemRLE),
    .io1_BranchJump_JrE(_mem2mem2_io1_BranchJump_JrE),
    .io1_Tlb_Control(_mem2mem2_io1_Tlb_Control),
    .io_en(_mem2mem2_io_en),
    .io_clr(_mem2mem2_io_clr),
    .io_WriteRegE(_mem2mem2_io_WriteRegE),
    .io_PhyAddrE(_mem2mem2_io_PhyAddrE),
    .io_HiLoOutE(_mem2mem2_io_HiLoOutE),
    .io_HiInE(_mem2mem2_io_HiInE),
    .io_LoInE(_mem2mem2_io_LoInE),
    .io_WriteCP0HiLoDataE(_mem2mem2_io_WriteCP0HiLoDataE),
    .io_BadVAddrE(_mem2mem2_io_BadVAddrE),
    .io_ExceptionTypeE(_mem2mem2_io_ExceptionTypeE),
    .io_RtE(_mem2mem2_io_RtE),
    .io_RegWriteM(_mem2mem2_io_RegWriteM),
    .io_MemToRegM(_mem2mem2_io_MemToRegM),
    .io_WriteRegM(_mem2mem2_io_WriteRegM),
    .io_LoadUnsignedM(_mem2mem2_io_LoadUnsignedM),
    .io_MemWidthM(_mem2mem2_io_MemWidthM),
    .io_PhyAddrM(_mem2mem2_io_PhyAddrM),
    .io_HiLoWriteM(_mem2mem2_io_HiLoWriteM),
    .io_HiLoOutM(_mem2mem2_io_HiLoOutM),
    .io_HiInM(_mem2mem2_io_HiInM),
    .io_LoInM(_mem2mem2_io_LoInM),
    .io_CP0WriteM(_mem2mem2_io_CP0WriteM),
    .io_WriteCP0AddrM(_mem2mem2_io_WriteCP0AddrM),
    .io_WriteCP0SelM(_mem2mem2_io_WriteCP0SelM),
    .io_WriteCP0HiLoDataM(_mem2mem2_io_WriteCP0HiLoDataM),
    .io_PCM(_mem2mem2_io_PCM),
    .io_InDelaySlotM(_mem2mem2_io_InDelaySlotM),
    .io_BadVAddrM(_mem2mem2_io_BadVAddrM),
    .io_ExceptionTypeM_Out(_mem2mem2_io_ExceptionTypeM_Out),
    .io_MemRLM(_mem2mem2_io_MemRLM),
    .io_RtM(_mem2mem2_io_RtM),
    .io_BranchJump_JrM(_mem2mem2_io_BranchJump_JrM),
    .io_Tlb_ControlM(_mem2mem2_io_Tlb_ControlM)
  );
  hilo _hilo ( // @[myCPU.scala 129:26]
    .clock(_hilo_clock),
    .reset(_hilo_reset),
    .io_we(_hilo_io_we),
    .io_hi_i(_hilo_io_hi_i),
    .io_lo_i(_hilo_io_lo_i),
    .io_hi_o(_hilo_io_hi_o),
    .io_lo_o(_hilo_io_lo_o)
  );
  id2ex _id2ex ( // @[myCPU.scala 130:26]
    .clock(_id2ex_clock),
    .reset(_id2ex_reset),
    .io1_RegWriteD(_id2ex_io1_RegWriteD),
    .io1_MemToRegD(_id2ex_io1_MemToRegD),
    .io1_MemWriteD(_id2ex_io1_MemWriteD),
    .io1_ALUCtrlD(_id2ex_io1_ALUCtrlD),
    .io1_ALUSrcD(_id2ex_io1_ALUSrcD),
    .io1_RegDstD(_id2ex_io1_RegDstD),
    .io1_LinkD(_id2ex_io1_LinkD),
    .io1_HiLoWriteD(_id2ex_io1_HiLoWriteD),
    .io1_HiLoToRegD(_id2ex_io1_HiLoToRegD),
    .io1_CP0WriteD(_id2ex_io1_CP0WriteD),
    .io1_CP0ToRegD(_id2ex_io1_CP0ToRegD),
    .io1_LoadUnsignedD(_id2ex_io1_LoadUnsignedD),
    .io1_MemWidthD(_id2ex_io1_MemWidthD),
    .io1_MemRLD(_id2ex_io1_MemRLD),
    .io2_RegWriteE(_id2ex_io2_RegWriteE),
    .io2_MemToRegE(_id2ex_io2_MemToRegE),
    .io2_MemWriteE(_id2ex_io2_MemWriteE),
    .io2_ALUCtrlE(_id2ex_io2_ALUCtrlE),
    .io2_ALUSrcE(_id2ex_io2_ALUSrcE),
    .io2_RegDstE(_id2ex_io2_RegDstE),
    .io2_LinkE(_id2ex_io2_LinkE),
    .io2_PCPlus8E(_id2ex_io2_PCPlus8E),
    .io2_LoadUnsignedE(_id2ex_io2_LoadUnsignedE),
    .io2_MemWidthE(_id2ex_io2_MemWidthE),
    .io2_HiLoWriteE(_id2ex_io2_HiLoWriteE),
    .io2_HiLoToRegE(_id2ex_io2_HiLoToRegE),
    .io2_CP0WriteE(_id2ex_io2_CP0WriteE),
    .io2_WriteCP0AddrE(_id2ex_io2_WriteCP0AddrE),
    .io2_WriteCP0SelE(_id2ex_io2_WriteCP0SelE),
    .io2_ReadCP0AddrE(_id2ex_io2_ReadCP0AddrE),
    .io2_ReadCP0SelE(_id2ex_io2_ReadCP0SelE),
    .io2_PCE(_id2ex_io2_PCE),
    .io2_InDelaySlotE(_id2ex_io2_InDelaySlotE),
    .io2_MemRLE(_id2ex_io2_MemRLE),
    .io2_BranchJump_JrE(_id2ex_io2_BranchJump_JrE),
    .io2_Tlb_Control(_id2ex_io2_Tlb_Control),
    .io_en(_id2ex_io_en),
    .io_clr(_id2ex_io_clr),
    .io_CP0ToRegE_Out(_id2ex_io_CP0ToRegE_Out),
    .io_RD1D(_id2ex_io_RD1D),
    .io_RD2D(_id2ex_io_RD2D),
    .io_RsD(_id2ex_io_RsD),
    .io_RtD(_id2ex_io_RtD),
    .io_RdD(_id2ex_io_RdD),
    .io_ImmD(_id2ex_io_ImmD),
    .io_PCPlus8D(_id2ex_io_PCPlus8D),
    .io_WriteCP0AddrD(_id2ex_io_WriteCP0AddrD),
    .io_WriteCP0SelD(_id2ex_io_WriteCP0SelD),
    .io_ReadCP0AddrD(_id2ex_io_ReadCP0AddrD),
    .io_ReadCP0SelD(_id2ex_io_ReadCP0SelD),
    .io_PCD(_id2ex_io_PCD),
    .io_InDelaySlotD(_id2ex_io_InDelaySlotD),
    .io_ExceptionTypeD(_id2ex_io_ExceptionTypeD),
    .io_BranchJump_JrD(_id2ex_io_BranchJump_JrD),
    .io_BadVaddrD(_id2ex_io_BadVaddrD),
    .io_Tlb_Control(_id2ex_io_Tlb_Control),
    .io_RD1E(_id2ex_io_RD1E),
    .io_RD2E(_id2ex_io_RD2E),
    .io_RsE(_id2ex_io_RsE),
    .io_RtE(_id2ex_io_RtE),
    .io_RdE(_id2ex_io_RdE),
    .io_ImmE(_id2ex_io_ImmE),
    .io_BadVaddrE(_id2ex_io_BadVaddrE),
    .io_ExceptionTypeE_Out(_id2ex_io_ExceptionTypeE_Out)
  );
  if2id _if2id ( // @[myCPU.scala 131:26]
    .clock(_if2id_clock),
    .reset(_if2id_reset),
    .io_en(_if2id_io_en),
    .io_clr(_if2id_io_clr),
    .io_InstrF(_if2id_io_InstrF),
    .io_PCPlus4F(_if2id_io_PCPlus4F),
    .io_PCPlus8F(_if2id_io_PCPlus8F),
    .io_PCF(_if2id_io_PCF),
    .io_ExceptionTypeF(_if2id_io_ExceptionTypeF),
    .io_NextDelaySlotD(_if2id_io_NextDelaySlotD),
    .io_InstrD(_if2id_io_InstrD),
    .io_PCPlus4D(_if2id_io_PCPlus4D),
    .io_PCPlus8D(_if2id_io_PCPlus8D),
    .io_InDelaySlotD(_if2id_io_InDelaySlotD),
    .io_PCD(_if2id_io_PCD),
    .io_ExceptionTypeD_Out(_if2id_io_ExceptionTypeD_Out)
  );
  mem2wb _mem22wb ( // @[myCPU.scala 133:27]
    .clock(_mem22wb_clock),
    .reset(_mem22wb_reset),
    .io_en(_mem22wb_io_en),
    .io_clr(_mem22wb_io_clr),
    .io_RegWriteM(_mem22wb_io_RegWriteM),
    .io_ResultM(_mem22wb_io_ResultM),
    .io_WriteRegM(_mem22wb_io_WriteRegM),
    .io_HiLoWriteM(_mem22wb_io_HiLoWriteM),
    .io_HiInM(_mem22wb_io_HiInM),
    .io_LoInM(_mem22wb_io_LoInM),
    .io_CP0WriteM(_mem22wb_io_CP0WriteM),
    .io_WriteCP0AddrM(_mem22wb_io_WriteCP0AddrM),
    .io_WriteCP0SelM(_mem22wb_io_WriteCP0SelM),
    .io_WriteCP0HiLoDataM(_mem22wb_io_WriteCP0HiLoDataM),
    .io_PCM(_mem22wb_io_PCM),
    .io_InDelaySlotM(_mem22wb_io_InDelaySlotM),
    .io_BadVAddrM(_mem22wb_io_BadVAddrM),
    .io_ExceptionTypeM(_mem22wb_io_ExceptionTypeM),
    .io_BranchJump_JrM(_mem22wb_io_BranchJump_JrM),
    .io_Tlb_ControlM(_mem22wb_io_Tlb_ControlM),
    .io_RegWriteW_Out(_mem22wb_io_RegWriteW_Out),
    .io_ResultW(_mem22wb_io_ResultW),
    .io_WriteRegW(_mem22wb_io_WriteRegW),
    .io_HiLoWriteW(_mem22wb_io_HiLoWriteW),
    .io_HiInW(_mem22wb_io_HiInW),
    .io_LoInW(_mem22wb_io_LoInW),
    .io_CP0WriteW(_mem22wb_io_CP0WriteW),
    .io_WriteCP0AddrW(_mem22wb_io_WriteCP0AddrW),
    .io_WriteCP0SelW(_mem22wb_io_WriteCP0SelW),
    .io_WriteCP0HiLoDataW(_mem22wb_io_WriteCP0HiLoDataW),
    .io_PCW(_mem22wb_io_PCW),
    .io_InDelaySlotW(_mem22wb_io_InDelaySlotW),
    .io_BadVAddrW(_mem22wb_io_BadVAddrW),
    .io_ExceptionTypeW_Out(_mem22wb_io_ExceptionTypeW_Out),
    .io_BranchJump_JrW(_mem22wb_io_BranchJump_JrW),
    .io_Tlb_ControlW(_mem22wb_io_Tlb_ControlW)
  );
  addr_cal _addr_cal ( // @[myCPU.scala 134:31]
    .io_d_vaddr(_addr_cal_io_d_vaddr),
    .io_d_width(_addr_cal_io_d_width),
    .io_d_memrl(_addr_cal_io_d_memrl),
    .io_d_paddr(_addr_cal_io_d_paddr),
    .io_d_cached(_addr_cal_io_d_cached),
    .io_d_unaligned(_addr_cal_io_d_unaligned)
  );
  muldiv _muldiv ( // @[myCPU.scala 135:26]
    .clock(_muldiv_clock),
    .reset(_muldiv_reset),
    .io_en(_muldiv_io_en),
    .io_ctrl(_muldiv_io_ctrl),
    .io_in1(_muldiv_io_in1),
    .io_in2(_muldiv_io_in2),
    .io_hi(_muldiv_io_hi),
    .io_lo(_muldiv_io_lo),
    .io_pending(_muldiv_io_pending)
  );
  regfile _regfile ( // @[myCPU.scala 137:26]
    .clock(_regfile_clock),
    .reset(_regfile_reset),
    .io_A1(_regfile_io_A1),
    .io_A2(_regfile_io_A2),
    .io_WE3(_regfile_io_WE3),
    .io_A3(_regfile_io_A3),
    .io_WD3(_regfile_io_WD3),
    .io_RD1(_regfile_io_RD1),
    .io_RD2(_regfile_io_RD2)
  );
  fifo fifo ( // @[myCPU.scala 139:29]
    .clock(fifo_clock),
    .reset(fifo_reset),
    .io_read_en(fifo_io_read_en),
    .io_write_en(fifo_io_write_en),
    .io_read_out_0(fifo_io_read_out_0),
    .io_write_in_0(fifo_io_write_in_0),
    .io_full(fifo_io_full),
    .io_empty(fifo_io_empty),
    .io_point_write_en(fifo_io_point_write_en),
    .io_point_flush(fifo_io_point_flush)
  );
  pc_detail stage_fec_1_pc_L ( // @[myCPU.scala 403:34]
    .clock(stage_fec_1_pc_L_clock),
    .reset(stage_fec_1_pc_L_reset),
    .io_stall(stage_fec_1_pc_L_io_stall),
    .io_flush(stage_fec_1_pc_L_io_flush),
    .io_in_pc_value_in(stage_fec_1_pc_L_io_in_pc_value_in),
    .io_out_pc_value_out(stage_fec_1_pc_L_io_out_pc_value_out)
  );
  pc_detail stage_fec_1_pc_M ( // @[myCPU.scala 404:34]
    .clock(stage_fec_1_pc_M_clock),
    .reset(stage_fec_1_pc_M_reset),
    .io_stall(stage_fec_1_pc_M_io_stall),
    .io_flush(stage_fec_1_pc_M_io_flush),
    .io_in_pc_value_in(stage_fec_1_pc_M_io_in_pc_value_in),
    .io_out_pc_value_out(stage_fec_1_pc_M_io_out_pc_value_out)
  );
  pc_detail stage_fec_1_pc_R ( // @[myCPU.scala 405:34]
    .clock(stage_fec_1_pc_R_clock),
    .reset(stage_fec_1_pc_R_reset),
    .io_stall(stage_fec_1_pc_R_io_stall),
    .io_flush(stage_fec_1_pc_R_io_flush),
    .io_in_pc_value_in(stage_fec_1_pc_R_io_in_pc_value_in),
    .io_out_pc_value_out(stage_fec_1_pc_R_io_out_pc_value_out)
  );
  branch_prediction_with_blockram branch_prediction_with_blockram ( // @[myCPU.scala 434:21]
    .clock(branch_prediction_with_blockram_clock),
    .reset(branch_prediction_with_blockram_reset),
    .io_pc(branch_prediction_with_blockram_io_pc),
    .io_write_pc(branch_prediction_with_blockram_io_write_pc),
    .io_aw_pht_ways_addr(branch_prediction_with_blockram_io_aw_pht_ways_addr),
    .io_aw_pht_addr(branch_prediction_with_blockram_io_aw_pht_addr),
    .io_aw_bht_addr(branch_prediction_with_blockram_io_aw_bht_addr),
    .io_aw_target_addr(branch_prediction_with_blockram_io_aw_target_addr),
    .io_btb_write(branch_prediction_with_blockram_io_btb_write),
    .io_bht_write(branch_prediction_with_blockram_io_bht_write),
    .io_pht_write(branch_prediction_with_blockram_io_pht_write),
    .io_bht_in(branch_prediction_with_blockram_io_bht_in),
    .io_pht_in(branch_prediction_with_blockram_io_pht_in),
    .io_out_L(branch_prediction_with_blockram_io_out_L),
    .io_pre_L(branch_prediction_with_blockram_io_pre_L),
    .io_bht_L(branch_prediction_with_blockram_io_bht_L),
    .io_btb_hit_0(branch_prediction_with_blockram_io_btb_hit_0),
    .io_pre_target_L(branch_prediction_with_blockram_io_pre_target_L),
    .io_stage2_stall(branch_prediction_with_blockram_io_stage2_stall),
    .io_stage2_flush(branch_prediction_with_blockram_io_stage2_flush),
    .io_pht_out(branch_prediction_with_blockram_io_pht_out),
    .io_lookup_data_0(branch_prediction_with_blockram_io_lookup_data_0)
  );
  pc_detail stage_fec_2_pc_L ( // @[myCPU.scala 503:34]
    .clock(stage_fec_2_pc_L_clock),
    .reset(stage_fec_2_pc_L_reset),
    .io_stall(stage_fec_2_pc_L_io_stall),
    .io_flush(stage_fec_2_pc_L_io_flush),
    .io_in_pc_value_in(stage_fec_2_pc_L_io_in_pc_value_in),
    .io_out_pc_value_out(stage_fec_2_pc_L_io_out_pc_value_out)
  );
  pc_detail stage_fec_2_pc_M ( // @[myCPU.scala 504:34]
    .clock(stage_fec_2_pc_M_clock),
    .reset(stage_fec_2_pc_M_reset),
    .io_stall(stage_fec_2_pc_M_io_stall),
    .io_flush(stage_fec_2_pc_M_io_flush),
    .io_in_pc_value_in(stage_fec_2_pc_M_io_in_pc_value_in),
    .io_out_pc_value_out(stage_fec_2_pc_M_io_out_pc_value_out)
  );
  pc_detail stage_fec_2_pc_R ( // @[myCPU.scala 505:34]
    .clock(stage_fec_2_pc_R_clock),
    .reset(stage_fec_2_pc_R_reset),
    .io_stall(stage_fec_2_pc_R_io_stall),
    .io_flush(stage_fec_2_pc_R_io_flush),
    .io_in_pc_value_in(stage_fec_2_pc_R_io_in_pc_value_in),
    .io_out_pc_value_out(stage_fec_2_pc_R_io_out_pc_value_out)
  );
  bru_detail id_bru_state ( // @[myCPU.scala 652:27]
    .clock(id_bru_state_clock),
    .reset(id_bru_state_reset),
    .io_stall(id_bru_state_io_stall),
    .io_flush(id_bru_state_io_flush),
    .io_in_pht(id_bru_state_io_in_pht),
    .io_in_bht(id_bru_state_io_in_bht),
    .io_in_hashcode(id_bru_state_io_in_hashcode),
    .io_in_target_pc(id_bru_state_io_in_target_pc),
    .io_in_lookup_data(id_bru_state_io_in_lookup_data),
    .io_in_pht_lookup_value(id_bru_state_io_in_pht_lookup_value),
    .io_out_pht(id_bru_state_io_out_pht),
    .io_out_bht(id_bru_state_io_out_bht),
    .io_out_hashcode(id_bru_state_io_out_hashcode),
    .io_out_target_pc(id_bru_state_io_out_target_pc),
    .io_out_lookup_data(id_bru_state_io_out_lookup_data),
    .io_out_pht_lookup_value(id_bru_state_io_out_pht_lookup_value)
  );
  bru_detail ex_bru_state ( // @[myCPU.scala 656:27]
    .clock(ex_bru_state_clock),
    .reset(ex_bru_state_reset),
    .io_stall(ex_bru_state_io_stall),
    .io_flush(ex_bru_state_io_flush),
    .io_in_pht(ex_bru_state_io_in_pht),
    .io_in_bht(ex_bru_state_io_in_bht),
    .io_in_hashcode(ex_bru_state_io_in_hashcode),
    .io_in_target_pc(ex_bru_state_io_in_target_pc),
    .io_in_lookup_data(ex_bru_state_io_in_lookup_data),
    .io_in_pht_lookup_value(ex_bru_state_io_in_pht_lookup_value),
    .io_out_pht(ex_bru_state_io_out_pht),
    .io_out_bht(ex_bru_state_io_out_bht),
    .io_out_hashcode(ex_bru_state_io_out_hashcode),
    .io_out_target_pc(ex_bru_state_io_out_target_pc),
    .io_out_lookup_data(ex_bru_state_io_out_lookup_data),
    .io_out_pht_lookup_value(ex_bru_state_io_out_pht_lookup_value)
  );
  bru_detail mem_bru_state ( // @[myCPU.scala 660:28]
    .clock(mem_bru_state_clock),
    .reset(mem_bru_state_reset),
    .io_stall(mem_bru_state_io_stall),
    .io_flush(mem_bru_state_io_flush),
    .io_in_pht(mem_bru_state_io_in_pht),
    .io_in_bht(mem_bru_state_io_in_bht),
    .io_in_hashcode(mem_bru_state_io_in_hashcode),
    .io_in_target_pc(mem_bru_state_io_in_target_pc),
    .io_in_lookup_data(mem_bru_state_io_in_lookup_data),
    .io_in_pht_lookup_value(mem_bru_state_io_in_pht_lookup_value),
    .io_out_pht(mem_bru_state_io_out_pht),
    .io_out_bht(mem_bru_state_io_out_bht),
    .io_out_hashcode(mem_bru_state_io_out_hashcode),
    .io_out_target_pc(mem_bru_state_io_out_target_pc),
    .io_out_lookup_data(mem_bru_state_io_out_lookup_data),
    .io_out_pht_lookup_value(mem_bru_state_io_out_pht_lookup_value)
  );
  bru_detail mem2_bru_state ( // @[myCPU.scala 664:29]
    .clock(mem2_bru_state_clock),
    .reset(mem2_bru_state_reset),
    .io_stall(mem2_bru_state_io_stall),
    .io_flush(mem2_bru_state_io_flush),
    .io_in_pht(mem2_bru_state_io_in_pht),
    .io_in_bht(mem2_bru_state_io_in_bht),
    .io_in_hashcode(mem2_bru_state_io_in_hashcode),
    .io_in_target_pc(mem2_bru_state_io_in_target_pc),
    .io_in_lookup_data(mem2_bru_state_io_in_lookup_data),
    .io_in_pht_lookup_value(mem2_bru_state_io_in_pht_lookup_value),
    .io_out_pht(mem2_bru_state_io_out_pht),
    .io_out_bht(mem2_bru_state_io_out_bht),
    .io_out_hashcode(mem2_bru_state_io_out_hashcode),
    .io_out_target_pc(mem2_bru_state_io_out_target_pc),
    .io_out_lookup_data(mem2_bru_state_io_out_lookup_data),
    .io_out_pht_lookup_value(mem2_bru_state_io_out_pht_lookup_value)
  );
  bru_detail wb_bru_state ( // @[myCPU.scala 668:27]
    .clock(wb_bru_state_clock),
    .reset(wb_bru_state_reset),
    .io_stall(wb_bru_state_io_stall),
    .io_flush(wb_bru_state_io_flush),
    .io_in_pht(wb_bru_state_io_in_pht),
    .io_in_bht(wb_bru_state_io_in_bht),
    .io_in_hashcode(wb_bru_state_io_in_hashcode),
    .io_in_target_pc(wb_bru_state_io_in_target_pc),
    .io_in_lookup_data(wb_bru_state_io_in_lookup_data),
    .io_in_pht_lookup_value(wb_bru_state_io_in_pht_lookup_value),
    .io_out_pht(wb_bru_state_io_out_pht),
    .io_out_bht(wb_bru_state_io_out_bht),
    .io_out_hashcode(wb_bru_state_io_out_hashcode),
    .io_out_target_pc(wb_bru_state_io_out_target_pc),
    .io_out_lookup_data(wb_bru_state_io_out_lookup_data),
    .io_out_pht_lookup_value(wb_bru_state_io_out_pht_lookup_value)
  );
  tlb_data_register tlb_data_register ( // @[myCPU.scala 971:30]
    .clock(tlb_data_register_clock),
    .reset(tlb_data_register_reset),
    .io_flush(tlb_data_register_io_flush),
    .io_stall(tlb_data_register_io_stall),
    .io_tlb_read_data_vaddr(tlb_data_register_io_tlb_read_data_vaddr),
    .io_tlb_read_data_asid(tlb_data_register_io_tlb_read_data_asid),
    .io_tlb_read_data_g(tlb_data_register_io_tlb_read_data_g),
    .io_tlb_read_data_paddr_0(tlb_data_register_io_tlb_read_data_paddr_0),
    .io_tlb_read_data_paddr_1(tlb_data_register_io_tlb_read_data_paddr_1),
    .io_tlb_read_data_c_0(tlb_data_register_io_tlb_read_data_c_0),
    .io_tlb_read_data_c_1(tlb_data_register_io_tlb_read_data_c_1),
    .io_tlb_read_data_d_0(tlb_data_register_io_tlb_read_data_d_0),
    .io_tlb_read_data_d_1(tlb_data_register_io_tlb_read_data_d_1),
    .io_tlb_read_data_v_0(tlb_data_register_io_tlb_read_data_v_0),
    .io_tlb_read_data_v_1(tlb_data_register_io_tlb_read_data_v_1),
    .io_tlb_write_data_vaddr(tlb_data_register_io_tlb_write_data_vaddr),
    .io_tlb_write_data_asid(tlb_data_register_io_tlb_write_data_asid),
    .io_tlb_write_data_g(tlb_data_register_io_tlb_write_data_g),
    .io_tlb_write_data_paddr_0(tlb_data_register_io_tlb_write_data_paddr_0),
    .io_tlb_write_data_paddr_1(tlb_data_register_io_tlb_write_data_paddr_1),
    .io_tlb_write_data_c_0(tlb_data_register_io_tlb_write_data_c_0),
    .io_tlb_write_data_c_1(tlb_data_register_io_tlb_write_data_c_1),
    .io_tlb_write_data_d_0(tlb_data_register_io_tlb_write_data_d_0),
    .io_tlb_write_data_d_1(tlb_data_register_io_tlb_write_data_d_1),
    .io_tlb_write_data_v_0(tlb_data_register_io_tlb_write_data_v_0),
    .io_tlb_write_data_v_1(tlb_data_register_io_tlb_write_data_v_1)
  );
  assign inst_cache = Pc_Next[31:29] == 3'h4; // @[macros.scala 420:55]
  assign inst_sram_en = stage2_stall; // @[myCPU.scala 366:17]
  assign inst_sram_addr = _stage_fec_2_branch_answer_T_7 ? _cp0_io_return_pc : _Pc_Next_T_3; // @[myCPU.scala 359:19]
  assign inst_ready_branch = fifo_io_point_write_en; // @[myCPU.scala 326:31 555:21]
  assign inst_buffer_empty = fifo_io_empty; // @[myCPU.scala 446:23]
  assign cp0_asid = _cp0_io_asid; // @[myCPU.scala 1165:14]
  assign stage2_flush = fifo_io_point_write_en & _stage_fec_2_data_valid_T | _stage_fec_2_branch_answer_T_7; // @[myCPU.scala 539:72]
  assign stage1_valid_flush = ready_to_branch & _access_stage1_sram_valid_T_1 & inst_write_en == 2'h0 ? 2'h2 : {{1'd0},
    _access_stage1_sram_valid_T_9}; // @[myCPU.scala 548:98 549:28]
  assign inst_ready_to_use = Pc_Next[1:0] == 2'h0; // @[myCPU.scala 367:39]
  assign inst_buffer_full = fifo_io_full; // @[myCPU.scala 556:22]
  assign data_sram_en = _dmemreq_io_req & ~_dmem_io_data_pending; // @[myCPU.scala 206:56]
  assign data_sram_wen = _dmemreq_io_wr; // @[myCPU.scala 212:13]
  assign data_size = _dmemreq_io_size; // @[myCPU.scala 1162:21]
  assign data_sram_addr = _dmemreq_io_addr; // @[myCPU.scala 208:15]
  assign data_sram_wdata = _dmemreq_io_wdata; // @[myCPU.scala 209:22]
  assign data_cache = commit_cache_reg & _addr_cal_io_d_cached; // @[myCPU.scala 1161:36]
  assign data_wstrb = _dmemreq_io_wstrb; // @[myCPU.scala 210:16]
  assign tlbp_search_vaddr = {resultE2M_Reg[31:13],13'h0}; // @[Cat.scala 31:58]
  assign tlbp_search_en = _ex2mem_io_Tlb_ControlM[2]; // @[myCPU.scala 984:45]
  assign tlb_read_index = resultE2M_Reg[3:0]; // @[myCPU.scala 978:37]
  assign tlb_write_index = ResultW[3:0]; // @[myCPU.scala 1127:32]
  assign debug_wb_pc = _mem22wb_io_PCW; // @[myCPU.scala 285:17]
  assign debug_wb_rf_wen = reg_pc == _mem22wb_io_PCW ? 4'h0 : _debug_wb_rf_wen_T_2; // @[myCPU.scala 286:27]
  assign debug_wb_rf_wnum = _regfile_io_A3; // @[myCPU.scala 287:22]
  assign debug_wb_rf_wdata = _regfile_io_WD3; // @[myCPU.scala 288:23]
  assign cp0_tlb_read_data_vaddr = _cp0_io_cp0_tlb_read_data_vaddr; // @[myCPU.scala 1177:23]
  assign cp0_tlb_read_data_asid = _cp0_io_cp0_tlb_read_data_asid; // @[myCPU.scala 1177:23]
  assign cp0_tlb_read_data_g = _cp0_io_cp0_tlb_read_data_g; // @[myCPU.scala 1177:23]
  assign cp0_tlb_read_data_paddr_0 = _cp0_io_cp0_tlb_read_data_paddr_0; // @[myCPU.scala 1177:23]
  assign cp0_tlb_read_data_paddr_1 = _cp0_io_cp0_tlb_read_data_paddr_1; // @[myCPU.scala 1177:23]
  assign cp0_tlb_read_data_c_0 = _cp0_io_cp0_tlb_read_data_c_0; // @[myCPU.scala 1177:23]
  assign cp0_tlb_read_data_c_1 = _cp0_io_cp0_tlb_read_data_c_1; // @[myCPU.scala 1177:23]
  assign cp0_tlb_read_data_d_0 = _cp0_io_cp0_tlb_read_data_d_0; // @[myCPU.scala 1177:23]
  assign cp0_tlb_read_data_d_1 = _cp0_io_cp0_tlb_read_data_d_1; // @[myCPU.scala 1177:23]
  assign cp0_tlb_read_data_v_0 = _cp0_io_cp0_tlb_read_data_v_0; // @[myCPU.scala 1177:23]
  assign cp0_tlb_read_data_v_1 = _cp0_io_cp0_tlb_read_data_v_1; // @[myCPU.scala 1177:23]
  assign tlb_write_en = _mem22wb_io_Tlb_ControlW[0]; // @[myCPU.scala 1126:45]
  assign _alu_io_ctrl = _id2ex_io2_ALUCtrlE; // @[myCPU.scala 848:18]
  assign _alu_io_in1 = _id2ex_io2_ALUSrcE[1] ? _Src1E_T_3 : RD1ForWardE; // @[myCPU.scala 842:20]
  assign _alu_io_in2 = _id2ex_io2_ALUSrcE[0] ? _id2ex_io_ImmE : RD2ForWardE; // @[myCPU.scala 843:20]
  assign _br_reset = ~resetn; // @[myCPU.scala 106:41]
  assign _br_io_rs = _cfu_io_ForwardAD[0] ? resultE2M_Reg : _BranchRsD_T_2; // @[myCPU.scala 739:20]
  assign _br_io_rt = _cfu_io_ForwardBD[0] ? resultE2M_Reg : _BranchRtD_T_2; // @[myCPU.scala 741:20]
  assign _br_io_branch = pre_decoder_branchdata; // @[myCPU.scala 748:19]
  assign _cfu_reset = ~resetn; // @[myCPU.scala 106:41]
  assign _cfu_io_Inst_Fifo_Empty = fifo_io_empty; // @[myCPU.scala 542:29]
  assign _cfu_io_dmem_calD = _cu_io1_dmem_addr_cal; // @[myCPU.scala 800:23]
  assign _cfu_io_BranchD_Flag = pre_decoder_branchD_flag; // @[myCPU.scala 1201:26]
  assign _cfu_io_JRD = pre_decoder_jr; // @[myCPU.scala 1197:25]
  assign _cfu_io_CanBranchD = ~(id_exception | ex_exception | mem_exception | mem2_exception | wb_exception); // @[myCPU.scala 1198:111]
  assign _cfu_io_DivPendingE = _muldiv_io_pending; // @[myCPU.scala 1202:33]
  assign _cfu_io_DataPendingM = _dmem_io_data_pending; // @[myCPU.scala 1204:33]
  assign _cfu_io_InException = _cp0_io_exception; // @[myCPU.scala 1184:25]
  assign _cfu_io_WriteRegE = 2'h3 == _id2ex_io2_RegDstE ? 5'h0 : _WriteRegE_T_3; // @[Mux.scala 81:58]
  assign _cfu_io_RegWriteE = _id2ex_io2_RegWriteE; // @[myCPU.scala 1210:33]
  assign _cfu_io_HiLoToRegE = _id2ex_io2_HiLoToRegE; // @[myCPU.scala 1211:33]
  assign _cfu_io_CP0ToRegE = _id2ex_io_ExceptionTypeE_Out == 32'h0 & _id2ex_io_CP0ToRegE_Out; // @[myCPU.scala 844:24]
  assign _cfu_io_WriteRegM = _ex2mem_io_WriteRegM; // @[myCPU.scala 1214:33]
  assign _cfu_io_MemToRegM = _ex2mem_io_MemToRegM; // @[myCPU.scala 1215:33]
  assign _cfu_io_RegWriteM = _ex2mem_io_RegWriteM; // @[myCPU.scala 1216:33]
  assign _cfu_io_HiLoWriteM = _ex2mem_io_HiLoWriteM; // @[myCPU.scala 1218:33]
  assign _cfu_io_CP0WriteM = _ex2mem_io_CP0WriteM; // @[myCPU.scala 1217:33]
  assign _cfu_io_WriteRegM2 = _mem2mem2_io_WriteRegM; // @[myCPU.scala 1240:25]
  assign _cfu_io_MemToRegM2 = _mem2mem2_io_MemToRegM; // @[myCPU.scala 1241:25]
  assign _cfu_io_RegWriteM2 = _mem2mem2_io_RegWriteM; // @[myCPU.scala 1242:25]
  assign _cfu_io_HiLoWriteM2 = _mem2mem2_io_HiLoWriteM; // @[myCPU.scala 1243:25]
  assign _cfu_io_CP0WriteM2 = _mem2mem2_io_CP0WriteM; // @[myCPU.scala 1237:24]
  assign _cfu_io_WriteRegW = _mem22wb_io_WriteRegW; // @[myCPU.scala 1228:33]
  assign _cfu_io_RegWriteW = wb_exception ? 1'h0 : _mem22wb_io_RegWriteW_Out; // @[myCPU.scala 1115:21]
  assign _cfu_io_HiLoWriteW = _mem22wb_io_HiLoWriteW; // @[myCPU.scala 1227:33]
  assign _cfu_io_CP0WriteW = _mem22wb_io_CP0WriteW; // @[myCPU.scala 1226:33]
  assign _cfu_io_ReadCP0AddrE = _id2ex_io2_ReadCP0AddrE; // @[myCPU.scala 1220:34]
  assign _cfu_io_ReadCP0SelE = _id2ex_io2_ReadCP0SelE; // @[myCPU.scala 1221:32]
  assign _cfu_io_WriteCP0AddrM = _ex2mem_io_WriteCP0AddrM; // @[myCPU.scala 1223:34]
  assign _cfu_io_WriteCP0SelM = _ex2mem_io_WriteCP0SelM; // @[myCPU.scala 1224:33]
  assign _cfu_io_WriteCP0AddrM2 = _mem2mem2_io_WriteCP0AddrM; // @[myCPU.scala 1238:28]
  assign _cfu_io_WriteCP0SelM2 = _mem2mem2_io_WriteCP0SelM; // @[myCPU.scala 1239:28]
  assign _cfu_io_RsD = _if2id_io_InstrD[25:21]; // @[myCPU.scala 182:27]
  assign _cfu_io_RtD = _if2id_io_InstrD[20:16]; // @[myCPU.scala 183:27]
  assign _cfu_io_RsE = _id2ex_io_RsE; // @[myCPU.scala 1233:33]
  assign _cfu_io_RtE = _id2ex_io_RtE; // @[myCPU.scala 1234:33]
  assign _cp0_clock = clk; // @[myCPU.scala 106:23]
  assign _cp0_reset = ~resetn; // @[myCPU.scala 106:41]
  assign _cp0_io_cp0_read_addr = _id2ex_io2_ReadCP0AddrE; // @[myCPU.scala 912:27]
  assign _cp0_io_cp0_read_sel = _id2ex_io2_ReadCP0SelE; // @[myCPU.scala 913:26]
  assign _cp0_io_cp0_write_addr = _mem22wb_io_WriteCP0AddrW; // @[myCPU.scala 914:28]
  assign _cp0_io_cp0_write_sel = _mem22wb_io_WriteCP0SelW; // @[myCPU.scala 915:27]
  assign _cp0_io_cp0_write_data = _mem22wb_io_WriteCP0HiLoDataW; // @[myCPU.scala 916:28]
  assign _cp0_io_cp0_write_en = CP0WriteW | tlb_exception_co0_writeW; // @[myCPU.scala 1171:47]
  assign _cp0_io_int_i = int_instanceW; // @[myCPU.scala 1168:19]
  assign _cp0_io_pc = _PCW_Reg_T ? _mem22wb_io_PCW : PCW_Reg; // @[myCPU.scala 1169:25]
  assign _cp0_io_mem_bad_vaddr = _mem22wb_io_BadVAddrW; // @[myCPU.scala 1170:27]
  assign _cp0_io_exception_type_i = _mem22wb_io_ExceptionTypeW_Out; // @[myCPU.scala 1172:30]
  assign _cp0_io_in_delayslot = _PCW_Reg_T ? _mem22wb_io_InDelaySlotW : slot_Reg; // @[myCPU.scala 1173:35]
  assign _cp0_io_in_branchjump_jr = _PCW_Reg_T ? _mem22wb_io_BranchJump_JrW : branchjump_Jr_Reg; // @[myCPU.scala 1174:37]
  assign _cp0_io_cp0_tlb_write_data_vaddr = tlb_data_register_io_tlb_read_data_vaddr; // @[myCPU.scala 1178:32]
  assign _cp0_io_cp0_tlb_write_data_asid = tlb_data_register_io_tlb_read_data_asid; // @[myCPU.scala 1178:32]
  assign _cp0_io_cp0_tlb_write_data_g = tlb_data_register_io_tlb_read_data_g; // @[myCPU.scala 1178:32]
  assign _cp0_io_cp0_tlb_write_data_paddr_0 = tlb_data_register_io_tlb_read_data_paddr_0; // @[myCPU.scala 1178:32]
  assign _cp0_io_cp0_tlb_write_data_paddr_1 = tlb_data_register_io_tlb_read_data_paddr_1; // @[myCPU.scala 1178:32]
  assign _cp0_io_cp0_tlb_write_data_c_0 = tlb_data_register_io_tlb_read_data_c_0; // @[myCPU.scala 1178:32]
  assign _cp0_io_cp0_tlb_write_data_c_1 = tlb_data_register_io_tlb_read_data_c_1; // @[myCPU.scala 1178:32]
  assign _cp0_io_cp0_tlb_write_data_d_0 = tlb_data_register_io_tlb_read_data_d_0; // @[myCPU.scala 1178:32]
  assign _cp0_io_cp0_tlb_write_data_d_1 = tlb_data_register_io_tlb_read_data_d_1; // @[myCPU.scala 1178:32]
  assign _cp0_io_cp0_tlb_write_data_v_0 = tlb_data_register_io_tlb_read_data_v_0; // @[myCPU.scala 1178:32]
  assign _cp0_io_cp0_tlb_write_data_v_1 = tlb_data_register_io_tlb_read_data_v_1; // @[myCPU.scala 1178:32]
  assign _cp0_io_cp0_tlb_write_en = _mem2mem2_io_Tlb_ControlM[1]; // @[myCPU.scala 1179:61]
  assign _cp0_io_cp0_index_tlb_write_able = _mem22wb_io_Tlb_ControlW[2]; // @[myCPU.scala 1180:65]
  assign _cu_reset = ~resetn; // @[myCPU.scala 106:41]
  assign _cu_io1_InstrD = _if2id_io_InstrD; // @[myCPU.scala 737:20]
  assign _dmem_io_data_ok = data_stage2_stall; // @[myCPU.scala 235:25]
  assign _dmem_io_rdata = data_sram_rdata; // @[myCPU.scala 236:25]
  assign _dmem_io_Physisc_Address = _mem2mem2_io_PhyAddrM; // @[myCPU.scala 244:30]
  assign _dmem_io_WIDTH = _mem2mem2_io_MemWidthM; // @[myCPU.scala 238:25]
  assign _dmem_io_SIGN = ~_mem2mem2_io_LoadUnsignedM; // @[myCPU.scala 239:22]
  assign _dmemreq_io_en = ex_exception | mem_exception | mem2_exception | wb_exception ? 1'h0 : __dmemreq_io_en_T_6; // @[myCPU.scala 862:26]
  assign _dmemreq_io_MemWriteE = _id2ex_io2_MemWriteE; // @[myCPU.scala 868:27]
  assign _dmemreq_io_MemToRegE = _id2ex_io2_MemToRegE; // @[myCPU.scala 865:27]
  assign _dmemreq_io_MemWidthE = _id2ex_io2_MemWidthE; // @[myCPU.scala 866:27]
  assign _dmemreq_io_VAddrE = _addr_cal_io_d_paddr; // @[myCPU.scala 1156:23]
  assign _dmemreq_io_WriteDataE = Forward_Lock2E ? RD2ForWardE_r : RD2ForWardE_p; // @[myCPU.scala 820:23]
  assign _dmemreq_io_memrl = _id2ex_io2_MemRLE; // @[myCPU.scala 872:23]
  assign _ex2mem_clock = clk; // @[myCPU.scala 106:23]
  assign _ex2mem_reset = ~resetn; // @[myCPU.scala 106:41]
  assign _ex2mem_io1_RegWriteE = _id2ex_io2_RegWriteE; // @[myCPU.scala 145:15]
  assign _ex2mem_io1_MemToRegE = _id2ex_io2_MemToRegE; // @[myCPU.scala 145:15]
  assign _ex2mem_io1_LoadUnsignedE = _id2ex_io2_LoadUnsignedE; // @[myCPU.scala 145:15]
  assign _ex2mem_io1_MemWidthE = _id2ex_io2_MemWidthE; // @[myCPU.scala 145:15]
  assign _ex2mem_io1_HiLoWriteE = _id2ex_io2_HiLoWriteE; // @[myCPU.scala 145:15]
  assign _ex2mem_io1_CP0WriteE = _id2ex_io2_CP0WriteE; // @[myCPU.scala 145:15]
  assign _ex2mem_io1_WriteCP0AddrE = _id2ex_io2_WriteCP0AddrE; // @[myCPU.scala 145:15]
  assign _ex2mem_io1_WriteCP0SelE = _id2ex_io2_WriteCP0SelE; // @[myCPU.scala 145:15]
  assign _ex2mem_io1_PCE = _id2ex_io2_PCE; // @[myCPU.scala 145:15]
  assign _ex2mem_io1_InDelaySlotE = _id2ex_io2_InDelaySlotE; // @[myCPU.scala 145:15]
  assign _ex2mem_io1_MemRLE = _id2ex_io2_MemRLE; // @[myCPU.scala 145:15]
  assign _ex2mem_io1_BranchJump_JrE = _id2ex_io2_BranchJump_JrE; // @[myCPU.scala 145:15]
  assign _ex2mem_io1_Tlb_Control = _id2ex_io2_Tlb_Control; // @[myCPU.scala 145:15]
  assign _ex2mem_io_en = _cfu_io_StallE; // @[myCPU.scala 191:30]
  assign _ex2mem_io_clr = _cfu_io_FlushM; // @[myCPU.scala 192:30]
  assign _ex2mem_io_WriteRegE = 2'h3 == _id2ex_io2_RegDstE ? 5'h0 : _WriteRegE_T_3; // @[Mux.scala 81:58]
  assign _ex2mem_io_PhyAddrE = _addr_cal_io_d_paddr; // @[myCPU.scala 907:27]
  assign _ex2mem_io_HiLoOutE = __ex2mem_io_HiLoOutE_T_14 | __ex2mem_io_HiLoOutE_T_15; // @[Mux.scala 27:73]
  assign _ex2mem_io_HiInE = _id2ex_io2_HiLoWriteE == 2'h2 ? WriteCP0HiLoDataE : _muldiv_io_hi; // @[myCPU.scala 857:20]
  assign _ex2mem_io_LoInE = _id2ex_io2_HiLoWriteE == 2'h1 ? WriteCP0HiLoDataE : _muldiv_io_lo; // @[myCPU.scala 858:20]
  assign _ex2mem_io_WriteCP0HiLoDataE = _id2ex_io2_HiLoWriteE != 2'h0 ? RD1ForWardE : _WriteCP0HiLoDataE_T_2; // @[myCPU.scala 840:32]
  assign _ex2mem_io_BadVAddrE = __dmemreq_io_en_T_3 & (_temp_exceptionE_T_2 | _temp_exceptionE_T_6) ?
    _addr_cal_io_d_vaddr : _BadVAddrE_T_9; // @[myCPU.scala 892:20]
  assign _ex2mem_io_ExceptionTypeE = _GEN_23 | temp_exceptionE; // @[myCPU.scala 896:127]
  assign _ex2mem_io_RtE = Forward_Lock2E ? RD2ForWardE_r : RD2ForWardE_p; // @[myCPU.scala 820:23]
  assign _mem2mem2_clock = clk; // @[myCPU.scala 106:23]
  assign _mem2mem2_reset = ~resetn; // @[myCPU.scala 106:41]
  assign _mem2mem2_io1_RegWriteE = _ex2mem_io_RegWriteM; // @[myCPU.scala 1014:30]
  assign _mem2mem2_io1_MemToRegE = _ex2mem_io_MemToRegM; // @[myCPU.scala 1015:30]
  assign _mem2mem2_io1_LoadUnsignedE = _ex2mem_io_LoadUnsignedM; // @[myCPU.scala 1019:30]
  assign _mem2mem2_io1_MemWidthE = _ex2mem_io_MemWidthM; // @[myCPU.scala 1020:30]
  assign _mem2mem2_io1_HiLoWriteE = _ex2mem_io_HiLoWriteM; // @[myCPU.scala 1021:30]
  assign _mem2mem2_io1_CP0WriteE = __mem2mem2_io_CP0WriteE_T_2 | __mem2mem2_io_WriteCP0HiLoDataE_T; // @[myCPU.scala 1023:91]
  assign _mem2mem2_io1_WriteCP0AddrE = __mem2mem2_io_WriteCP0HiLoDataE_T | inst_tlb_exceptionM ? 5'ha :
    _ex2mem_io_WriteCP0AddrM; // @[myCPU.scala 1024:36]
  assign _mem2mem2_io1_WriteCP0SelE = __mem2mem2_io1_WriteCP0AddrE_T_1 ? 3'h0 : _ex2mem_io_WriteCP0SelM; // @[myCPU.scala 1025:36]
  assign _mem2mem2_io1_PCE = _ex2mem_io_PCM; // @[myCPU.scala 1026:30]
  assign _mem2mem2_io1_InDelaySlotE = _ex2mem_io_InDelaySlotM; // @[myCPU.scala 1027:30]
  assign _mem2mem2_io1_MemRLE = _ex2mem_io_MemRLM; // @[myCPU.scala 1028:30]
  assign _mem2mem2_io1_BranchJump_JrE = _ex2mem_io_BranchJump_JrM; // @[myCPU.scala 1029:30]
  assign _mem2mem2_io1_Tlb_Control = _ex2mem_io_Tlb_ControlM; // @[myCPU.scala 1039:27]
  assign _mem2mem2_io_en = _cfu_io_StallM2; // @[myCPU.scala 1059:20]
  assign _mem2mem2_io_clr = _cfu_io_FlushM2; // @[myCPU.scala 1058:20]
  assign _mem2mem2_io_WriteRegE = _ex2mem_io_WriteRegM; // @[myCPU.scala 998:24]
  assign _mem2mem2_io_PhyAddrE = _ex2mem_io_PhyAddrM; // @[myCPU.scala 999:23]
  assign _mem2mem2_io_HiLoOutE = _ex2mem_io_HiLoOutM; // @[myCPU.scala 1054:30]
  assign _mem2mem2_io_HiInE = _ex2mem_io_HiInM; // @[myCPU.scala 1000:20]
  assign _mem2mem2_io_LoInE = _ex2mem_io_LoInM; // @[myCPU.scala 1001:20]
  assign _mem2mem2_io_WriteCP0HiLoDataE = __mem2mem2_io_WriteCP0HiLoDataE_T ? __mem2mem2_io_WriteCP0HiLoDataE_T_2 :
    __mem2mem2_io_WriteCP0HiLoDataE_T_7; // @[Mux.scala 101:16]
  assign _mem2mem2_io_BadVAddrE = __mem2mem2_io_WriteCP0HiLoDataE_T ? _ex2mem_io_PhyAddrM : __mem2mem2_io_BadVAddrE_T_9; // @[myCPU.scala 1049:36]
  assign _mem2mem2_io_ExceptionTypeE = mem_exception ? _ex2mem_io_ExceptionTypeM_Out : {{24'd0}, _ExceptionM_T_11}; // @[myCPU.scala 992:21]
  assign _mem2mem2_io_RtE = _ex2mem_io_RtM; // @[myCPU.scala 1012:18]
  assign _hilo_clock = clk; // @[myCPU.scala 106:23]
  assign _hilo_reset = ~resetn; // @[myCPU.scala 106:41]
  assign _hilo_io_we = wb_exception ? 2'h0 : _mem22wb_io_HiLoWriteW; // @[myCPU.scala 1116:25]
  assign _hilo_io_hi_i = _mem22wb_io_HiInW; // @[myCPU.scala 918:19]
  assign _hilo_io_lo_i = _mem22wb_io_LoInW; // @[myCPU.scala 919:19]
  assign _id2ex_clock = clk; // @[myCPU.scala 106:23]
  assign _id2ex_reset = ~resetn; // @[myCPU.scala 106:41]
  assign _id2ex_io1_RegWriteD = _cu_io_RegWriteD; // @[myCPU.scala 144:15]
  assign _id2ex_io1_MemToRegD = _cu_io_MemToRegD; // @[myCPU.scala 144:15]
  assign _id2ex_io1_MemWriteD = _cu_io_MemWriteD; // @[myCPU.scala 144:15]
  assign _id2ex_io1_ALUCtrlD = _cu_io_ALUCtrlD; // @[myCPU.scala 144:15]
  assign _id2ex_io1_ALUSrcD = _cu_io_ALUSrcD; // @[myCPU.scala 144:15]
  assign _id2ex_io1_RegDstD = _cu_io_RegDstD; // @[myCPU.scala 144:15]
  assign _id2ex_io1_LinkD = _cu_io_LinkD; // @[myCPU.scala 144:15]
  assign _id2ex_io1_HiLoWriteD = _cu_io_HiLoWriteD; // @[myCPU.scala 144:15]
  assign _id2ex_io1_HiLoToRegD = _cu_io_HiLoToRegD; // @[myCPU.scala 144:15]
  assign _id2ex_io1_CP0WriteD = _cu_io_CP0WriteD; // @[myCPU.scala 144:15]
  assign _id2ex_io1_CP0ToRegD = _cu_io_CP0ToRegD; // @[myCPU.scala 144:15]
  assign _id2ex_io1_LoadUnsignedD = _cu_io_LoadUnsignedD; // @[myCPU.scala 144:15]
  assign _id2ex_io1_MemWidthD = _cu_io_MemWidthD; // @[myCPU.scala 144:15]
  assign _id2ex_io1_MemRLD = _cu_io_MemRLD; // @[myCPU.scala 144:15]
  assign _id2ex_io_en = _cfu_io_StallD; // @[myCPU.scala 172:29]
  assign _id2ex_io_clr = _cfu_io_FlushE; // @[myCPU.scala 173:29]
  assign _id2ex_io_RD1D = _cfu_io_ForwardAD[0] ? resultE2M_Reg : _BranchRsD_T_2; // @[myCPU.scala 777:25]
  assign _id2ex_io_RD2D = _cfu_io_ForwardBD[0] ? resultE2M_Reg : _BranchRtD_T_2; // @[myCPU.scala 778:25]
  assign _id2ex_io_RsD = _if2id_io_InstrD[25:21]; // @[myCPU.scala 182:27]
  assign _id2ex_io_RtD = _if2id_io_InstrD[20:16]; // @[myCPU.scala 183:27]
  assign _id2ex_io_RdD = _if2id_io_InstrD[15:11]; // @[myCPU.scala 184:27]
  assign _id2ex_io_ImmD = _cu_io_ImmUnsigned ? {{15'd0}, _ImmD_T_3} : _ImmD_T_23; // @[myCPU.scala 185:24]
  assign _id2ex_io_PCPlus8D = _if2id_io_PCPlus8D; // @[myCPU.scala 789:29]
  assign _id2ex_io_WriteCP0AddrD = _cu_io1_Tlb_Control[2] ? 5'h0 : RdD; // @[myCPU.scala 779:35]
  assign _id2ex_io_WriteCP0SelD = _cu_io1_Tlb_Control[2] ? 3'h0 : Write_WriteCP0Sel0; // @[myCPU.scala 780:35]
  assign _id2ex_io_ReadCP0AddrD = __if2id_io_InstrF_T_5 ? 5'he : __id2ex_io_ReadCP0AddrD_T_7; // @[Mux.scala 101:16]
  assign _id2ex_io_ReadCP0SelD = __if2id_io_InstrF_T_5 | _cu_io1_Tlb_Control[2] | _cu_io1_Tlb_Control[1] |
    _cu_io1_Tlb_Control[0] ? 3'h0 : Write_WriteCP0Sel0; // @[myCPU.scala 788:35]
  assign _id2ex_io_PCD = _if2id_io_PCD; // @[myCPU.scala 791:28]
  assign _id2ex_io_InDelaySlotD = _if2id_io_InDelaySlotD & _if2id_io_PCD[1:0] == 2'h0; // @[myCPU.scala 790:61]
  assign _id2ex_io_ExceptionTypeD = __id2ex_io_ExceptionTypeD_T != 6'h0 & _cp0_io_Int_able ? 32'h1 :
    __id2ex_io_ExceptionTypeD_T_16; // @[myCPU.scala 767:37]
  assign _id2ex_io_BranchJump_JrD = {1'h0,_T_54}; // @[Cat.scala 31:58]
  assign _id2ex_io_BadVaddrD = _if2id_io_PCD; // @[myCPU.scala 794:28]
  assign _id2ex_io_Tlb_Control = _cu_io1_Tlb_Control; // @[myCPU.scala 795:28]
  assign _if2id_clock = clk; // @[myCPU.scala 106:23]
  assign _if2id_reset = ~resetn; // @[myCPU.scala 106:41]
  assign _if2id_io_en = _cfu_io_StallD; // @[myCPU.scala 580:30]
  assign _if2id_io_clr = _cfu_io_FlushD; // @[myCPU.scala 581:30]
  assign _if2id_io_InstrF = _cu_io1_BadInstrD | _cu_io1_SysCallD | _cu_io1_BreakD | __if2id_io_InstrF_T_5 ? 32'h0 :
    fifo_io_read_out_0[63:32]; // @[myCPU.scala 584:33]
  assign _if2id_io_PCPlus4F = _if2id_io_PCF + 32'h4; // @[myCPU.scala 578:48]
  assign _if2id_io_PCPlus8F = _if2id_io_PCF + 32'h8; // @[myCPU.scala 579:48]
  assign _if2id_io_PCF = fifo_io_read_out_0[31:0]; // @[myCPU.scala 577:57]
  assign _if2id_io_ExceptionTypeF = fifo_io_read_out_0[135:134]; // @[myCPU.scala 582:56]
  assign _if2id_io_NextDelaySlotD = _T_54 | InDelaySlotF; // @[myCPU.scala 587:94]
  assign _mem22wb_clock = clk; // @[myCPU.scala 106:23]
  assign _mem22wb_reset = ~resetn; // @[myCPU.scala 106:41]
  assign _mem22wb_io_en = _cfu_io_StallW; // @[myCPU.scala 248:31]
  assign _mem22wb_io_clr = _cfu_io_FlushW; // @[myCPU.scala 249:31]
  assign _mem22wb_io_RegWriteM = _mem2mem2_io_RegWriteM; // @[myCPU.scala 251:38]
  assign _mem22wb_io_ResultM = _Forward_Lock1E_T_1 ? Mem_withRL_Data : ResultM2_Reg; // @[myCPU.scala 1069:25]
  assign _mem22wb_io_WriteRegM = _mem2mem2_io_WriteRegM; // @[myCPU.scala 253:38]
  assign _mem22wb_io_HiLoWriteM = _mem2mem2_io_HiLoWriteM; // @[myCPU.scala 263:38]
  assign _mem22wb_io_HiInM = _mem2mem2_io_HiInM; // @[myCPU.scala 254:38]
  assign _mem22wb_io_LoInM = _mem2mem2_io_LoInM; // @[myCPU.scala 255:38]
  assign _mem22wb_io_CP0WriteM = _mem2mem2_io_CP0WriteM; // @[myCPU.scala 259:38]
  assign _mem22wb_io_WriteCP0AddrM = _mem2mem2_io_WriteCP0AddrM; // @[myCPU.scala 260:38]
  assign _mem22wb_io_WriteCP0SelM = _mem2mem2_io_WriteCP0SelM; // @[myCPU.scala 261:38]
  assign _mem22wb_io_WriteCP0HiLoDataM = _mem2mem2_io_WriteCP0HiLoDataM; // @[myCPU.scala 262:38]
  assign _mem22wb_io_PCM = _mem2mem2_io_PCM; // @[myCPU.scala 258:38]
  assign _mem22wb_io_InDelaySlotM = _mem2mem2_io_InDelaySlotM; // @[myCPU.scala 256:38]
  assign _mem22wb_io_BadVAddrM = _mem2mem2_io_BadVAddrM; // @[myCPU.scala 1093:30]
  assign _mem22wb_io_ExceptionTypeM = _mem2mem2_io_ExceptionTypeM_Out; // @[myCPU.scala 1085:33]
  assign _mem22wb_io_BranchJump_JrM = _mem2mem2_io_BranchJump_JrM; // @[myCPU.scala 1089:33]
  assign _mem22wb_io_Tlb_ControlM = _mem2mem2_io_Tlb_ControlM; // @[myCPU.scala 264:38]
  assign _addr_cal_io_d_vaddr = _id2ex_io_ImmE + _id2ex_io_RD1E; // @[myCPU.scala 1154:44]
  assign _addr_cal_io_d_width = _id2ex_io2_MemWidthE; // @[myCPU.scala 1153:26]
  assign _addr_cal_io_d_memrl = _id2ex_io2_MemRLE; // @[myCPU.scala 1157:25]
  assign _muldiv_clock = clk; // @[myCPU.scala 106:23]
  assign _muldiv_reset = ~resetn; // @[myCPU.scala 106:41]
  assign _muldiv_io_en = ~ex_exception; // @[myCPU.scala 850:22]
  assign _muldiv_io_ctrl = {_muldiv_io_ctrl_hi,_id2ex_io2_ALUCtrlE[6:5]}; // @[Cat.scala 31:58]
  assign _muldiv_io_in1 = _id2ex_io2_ALUSrcE[1] ? _Src1E_T_3 : RD1ForWardE; // @[myCPU.scala 842:20]
  assign _muldiv_io_in2 = _id2ex_io2_ALUSrcE[0] ? _id2ex_io_ImmE : RD2ForWardE; // @[myCPU.scala 843:20]
  assign _regfile_clock = clk; // @[myCPU.scala 106:23]
  assign _regfile_reset = ~resetn; // @[myCPU.scala 106:41]
  assign _regfile_io_A1 = _if2id_io_InstrD[25:21]; // @[myCPU.scala 735:29]
  assign _regfile_io_A2 = _if2id_io_InstrD[20:16]; // @[myCPU.scala 736:29]
  assign _regfile_io_WE3 = wb_exception ? 1'h0 : _mem22wb_io_RegWriteW_Out; // @[myCPU.scala 1115:21]
  assign _regfile_io_A3 = _mem22wb_io_WriteRegW; // @[myCPU.scala 1121:21]
  assign _regfile_io_WD3 = _mem22wb_io_ResultW; // @[myCPU.scala 1114:15 270:26]
  assign fifo_clock = clk; // @[myCPU.scala 106:23]
  assign fifo_reset = ~resetn; // @[myCPU.scala 106:41]
  assign fifo_io_read_en = {{1'd0}, _T_35}; // @[myCPU.scala 535:29]
  assign fifo_io_write_en = inst_write_en; // @[myCPU.scala 531:35]
  assign fifo_io_write_in_0 = {hi,lo}; // @[Cat.scala 31:58]
  assign fifo_io_point_write_en = _PCSrcD_T_1 & ((pre_decoder_jump | _PCSrcD_T_3) != id_true_branch_state |
    target_addr_error); // @[myCPU.scala 699:57]
  assign fifo_io_point_flush = _cp0_io_exception; // @[myCPU.scala 536:29]
  assign stage_fec_1_pc_L_clock = clk; // @[myCPU.scala 106:23]
  assign stage_fec_1_pc_L_reset = ~resetn; // @[myCPU.scala 106:41]
  assign stage_fec_1_pc_L_io_stall = stage2_stall; // @[myCPU.scala 426:31]
  assign stage_fec_1_pc_L_io_flush = _stage_fec_2_branch_answer_T_7 & ~stage2_stall; // @[myCPU.scala 384:54]
  assign stage_fec_1_pc_L_io_in_pc_value_in = _stage_fec_2_branch_answer_T_7 ? _cp0_io_return_pc : _Pc_Next_T_3; // @[myCPU.scala 359:19]
  assign stage_fec_1_pc_M_clock = clk; // @[myCPU.scala 106:23]
  assign stage_fec_1_pc_M_reset = ~resetn; // @[myCPU.scala 106:41]
  assign stage_fec_1_pc_M_io_stall = stage2_stall; // @[myCPU.scala 427:31]
  assign stage_fec_1_pc_M_io_flush = _stage_fec_2_branch_answer_T_7 & ~stage2_stall; // @[myCPU.scala 384:54]
  assign stage_fec_1_pc_M_io_in_pc_value_in = _stage_fec_2_branch_answer_T_7 ? _cp0_io_return_pc : _Pc_Next_T_3; // @[myCPU.scala 359:19]
  assign stage_fec_1_pc_R_clock = clk; // @[myCPU.scala 106:23]
  assign stage_fec_1_pc_R_reset = ~resetn; // @[myCPU.scala 106:41]
  assign stage_fec_1_pc_R_io_stall = stage2_stall; // @[myCPU.scala 428:31]
  assign stage_fec_1_pc_R_io_flush = _stage_fec_2_branch_answer_T_7 & ~stage2_stall; // @[myCPU.scala 384:54]
  assign stage_fec_1_pc_R_io_in_pc_value_in = _stage_fec_2_branch_answer_T_7 ? _cp0_io_return_pc : _Pc_Next_T_3; // @[myCPU.scala 359:19]
  assign branch_prediction_with_blockram_clock = clk; // @[myCPU.scala 106:23]
  assign branch_prediction_with_blockram_reset = ~resetn; // @[myCPU.scala 106:41]
  assign branch_prediction_with_blockram_io_pc = stage_fec_1_pc_L_io_out_pc_value_out; // @[myCPU.scala 435:12]
  assign branch_prediction_with_blockram_io_write_pc = _mem22wb_io_PCW; // @[myCPU.scala 1139:17]
  assign branch_prediction_with_blockram_io_aw_pht_ways_addr = wb_bru_state_io_out_hashcode; // @[myCPU.scala 1138:25]
  assign branch_prediction_with_blockram_io_aw_pht_addr = wb_bru_state_io_out_lookup_data; // @[myCPU.scala 1136:20]
  assign branch_prediction_with_blockram_io_aw_bht_addr = _mem22wb_io_PCW[10:4]; // @[myCPU.scala 1135:38]
  assign branch_prediction_with_blockram_io_aw_target_addr = wb_bru_state_io_out_target_pc; // @[myCPU.scala 1137:23]
  assign branch_prediction_with_blockram_io_btb_write = branch_prediction_with_blockram_io_bht_write; // @[myCPU.scala 1134:18]
  assign branch_prediction_with_blockram_io_bht_write = _mem22wb_io_BranchJump_JrW[0]; // @[myCPU.scala 1132:47]
  assign branch_prediction_with_blockram_io_pht_write = branch_prediction_with_blockram_io_bht_write; // @[myCPU.scala 1133:18]
  assign branch_prediction_with_blockram_io_bht_in = wb_bru_state_io_out_bht; // @[myCPU.scala 1130:15]
  assign branch_prediction_with_blockram_io_pht_in = wb_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 1131:15]
  assign branch_prediction_with_blockram_io_stage2_stall = stage2_stall; // @[myCPU.scala 458:22]
  assign branch_prediction_with_blockram_io_stage2_flush = stage2_flush; // @[myCPU.scala 457:22]
  assign stage_fec_2_pc_L_clock = clk; // @[myCPU.scala 106:23]
  assign stage_fec_2_pc_L_reset = ~resetn; // @[myCPU.scala 106:41]
  assign stage_fec_2_pc_L_io_stall = stage2_stall; // @[myCPU.scala 527:31]
  assign stage_fec_2_pc_L_io_flush = stage2_flush; // @[myCPU.scala 523:31]
  assign stage_fec_2_pc_L_io_in_pc_value_in = stage_fec_1_pc_L_io_out_pc_value_out; // @[myCPU.scala 514:40]
  assign stage_fec_2_pc_M_clock = clk; // @[myCPU.scala 106:23]
  assign stage_fec_2_pc_M_reset = ~resetn; // @[myCPU.scala 106:41]
  assign stage_fec_2_pc_M_io_stall = stage2_stall; // @[myCPU.scala 528:31]
  assign stage_fec_2_pc_M_io_flush = stage2_flush; // @[myCPU.scala 524:31]
  assign stage_fec_2_pc_M_io_in_pc_value_in = stage_fec_1_pc_M_io_out_pc_value_out; // @[myCPU.scala 517:40]
  assign stage_fec_2_pc_R_clock = clk; // @[myCPU.scala 106:23]
  assign stage_fec_2_pc_R_reset = ~resetn; // @[myCPU.scala 106:41]
  assign stage_fec_2_pc_R_io_stall = stage2_stall; // @[myCPU.scala 529:31]
  assign stage_fec_2_pc_R_io_flush = stage2_flush; // @[myCPU.scala 525:31]
  assign stage_fec_2_pc_R_io_in_pc_value_in = stage_fec_1_pc_R_io_out_pc_value_out; // @[myCPU.scala 520:40]
  assign id_bru_state_clock = clk; // @[myCPU.scala 106:23]
  assign id_bru_state_reset = ~resetn; // @[myCPU.scala 106:41]
  assign id_bru_state_io_stall = _cfu_io_StallD; // @[myCPU.scala 654:23]
  assign id_bru_state_io_flush = _cfu_io_FlushD; // @[myCPU.scala 653:23]
  assign id_bru_state_io_in_pht = fifo_io_read_out_0[108:107]; // @[myCPU.scala 685:54]
  assign id_bru_state_io_in_bht = fifo_io_read_out_0[115:109]; // @[myCPU.scala 686:54]
  assign id_bru_state_io_in_hashcode = fifo_io_read_out_0[74:71]; // @[myCPU.scala 683:59]
  assign id_bru_state_io_in_target_pc = fifo_io_read_out_0[106:75]; // @[myCPU.scala 684:60]
  assign id_bru_state_io_in_lookup_data = fifo_io_read_out_0[70:64]; // @[myCPU.scala 682:62]
  assign id_bru_state_io_in_pht_lookup_value = fifo_io_read_out_0[124:117]; // @[myCPU.scala 687:67]
  assign ex_bru_state_clock = clk; // @[myCPU.scala 106:23]
  assign ex_bru_state_reset = ~resetn; // @[myCPU.scala 106:41]
  assign ex_bru_state_io_stall = _cfu_io_StallE; // @[myCPU.scala 658:23]
  assign ex_bru_state_io_flush = _cfu_io_FlushE; // @[myCPU.scala 657:23]
  assign ex_bru_state_io_in_pht = id_bru_state_io_out_pht; // @[myCPU.scala 715:28]
  assign ex_bru_state_io_in_bht = id_bru_state_io_out_bht; // @[myCPU.scala 714:28]
  assign ex_bru_state_io_in_hashcode = id_bru_state_io_out_hashcode; // @[myCPU.scala 716:33]
  assign ex_bru_state_io_in_target_pc = pre_decoder_branchD_flag ? PCBranchD : _Pc_targetD_T_2; // @[Mux.scala 101:16]
  assign ex_bru_state_io_in_lookup_data = id_bru_state_io_out_lookup_data; // @[myCPU.scala 717:36]
  assign ex_bru_state_io_in_pht_lookup_value = id_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 718:41]
  assign mem_bru_state_clock = clk; // @[myCPU.scala 106:23]
  assign mem_bru_state_reset = ~resetn; // @[myCPU.scala 106:41]
  assign mem_bru_state_io_stall = _cfu_io_StallM; // @[myCPU.scala 662:24]
  assign mem_bru_state_io_flush = _cfu_io_FlushM; // @[myCPU.scala 661:24]
  assign mem_bru_state_io_in_pht = 2'h2 == ex_bru_state_io_out_pht ? _pht_tobeE_T_3 : _pht_tobeE_T_7; // @[Mux.scala 81:58]
  assign mem_bru_state_io_in_bht = {ex_bru_state_io_out_bht[5:0],true_branch_stateE}; // @[Cat.scala 31:58]
  assign mem_bru_state_io_in_hashcode = ex_bru_state_io_out_hashcode; // @[myCPU.scala 673:22]
  assign mem_bru_state_io_in_target_pc = ex_bru_state_io_out_target_pc; // @[myCPU.scala 673:22]
  assign mem_bru_state_io_in_lookup_data = ex_bru_state_io_out_lookup_data; // @[myCPU.scala 673:22]
  assign mem_bru_state_io_in_pht_lookup_value = 2'h3 == ex_bru_state_io_out_lookup_data[1:0] ?
    _pht_lookup_value_tobeE_T_10 : _pht_lookup_value_tobeE_T_14; // @[Mux.scala 81:58]
  assign mem2_bru_state_clock = clk; // @[myCPU.scala 106:23]
  assign mem2_bru_state_reset = ~resetn; // @[myCPU.scala 106:41]
  assign mem2_bru_state_io_stall = _cfu_io_StallM2; // @[myCPU.scala 666:25]
  assign mem2_bru_state_io_flush = _cfu_io_FlushM2; // @[myCPU.scala 665:25]
  assign mem2_bru_state_io_in_pht = mem_bru_state_io_out_pht; // @[myCPU.scala 674:22]
  assign mem2_bru_state_io_in_bht = mem_bru_state_io_out_bht; // @[myCPU.scala 674:22]
  assign mem2_bru_state_io_in_hashcode = mem_bru_state_io_out_hashcode; // @[myCPU.scala 674:22]
  assign mem2_bru_state_io_in_target_pc = mem_bru_state_io_out_target_pc; // @[myCPU.scala 674:22]
  assign mem2_bru_state_io_in_lookup_data = mem_bru_state_io_out_lookup_data; // @[myCPU.scala 674:22]
  assign mem2_bru_state_io_in_pht_lookup_value = mem_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 674:22]
  assign wb_bru_state_clock = clk; // @[myCPU.scala 106:23]
  assign wb_bru_state_reset = ~resetn; // @[myCPU.scala 106:41]
  assign wb_bru_state_io_stall = _cfu_io_StallW; // @[myCPU.scala 670:23]
  assign wb_bru_state_io_flush = _cfu_io_FlushW; // @[myCPU.scala 669:23]
  assign wb_bru_state_io_in_pht = mem2_bru_state_io_out_pht; // @[myCPU.scala 675:22]
  assign wb_bru_state_io_in_bht = mem2_bru_state_io_out_bht; // @[myCPU.scala 675:22]
  assign wb_bru_state_io_in_hashcode = mem2_bru_state_io_out_hashcode; // @[myCPU.scala 675:22]
  assign wb_bru_state_io_in_target_pc = mem2_bru_state_io_out_target_pc; // @[myCPU.scala 675:22]
  assign wb_bru_state_io_in_lookup_data = mem2_bru_state_io_out_lookup_data; // @[myCPU.scala 675:22]
  assign wb_bru_state_io_in_pht_lookup_value = mem2_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 675:22]
  assign tlb_data_register_clock = clk; // @[myCPU.scala 106:23]
  assign tlb_data_register_reset = ~resetn; // @[myCPU.scala 106:41]
  assign tlb_data_register_io_flush = _cfu_io_FlushM2; // @[myCPU.scala 972:23]
  assign tlb_data_register_io_stall = _cfu_io_StallM2; // @[myCPU.scala 973:23]
  assign tlb_data_register_io_tlb_write_data_vaddr = cp0_tlb_write_data_vaddr; // @[myCPU.scala 974:32]
  assign tlb_data_register_io_tlb_write_data_asid = cp0_tlb_write_data_asid; // @[myCPU.scala 974:32]
  assign tlb_data_register_io_tlb_write_data_g = cp0_tlb_write_data_g; // @[myCPU.scala 974:32]
  assign tlb_data_register_io_tlb_write_data_paddr_0 = cp0_tlb_write_data_paddr_0; // @[myCPU.scala 974:32]
  assign tlb_data_register_io_tlb_write_data_paddr_1 = cp0_tlb_write_data_paddr_1; // @[myCPU.scala 974:32]
  assign tlb_data_register_io_tlb_write_data_c_0 = cp0_tlb_write_data_c_0; // @[myCPU.scala 974:32]
  assign tlb_data_register_io_tlb_write_data_c_1 = cp0_tlb_write_data_c_1; // @[myCPU.scala 974:32]
  assign tlb_data_register_io_tlb_write_data_d_0 = cp0_tlb_write_data_d_0; // @[myCPU.scala 974:32]
  assign tlb_data_register_io_tlb_write_data_d_1 = cp0_tlb_write_data_d_1; // @[myCPU.scala 974:32]
  assign tlb_data_register_io_tlb_write_data_v_0 = cp0_tlb_write_data_v_0; // @[myCPU.scala 974:32]
  assign tlb_data_register_io_tlb_write_data_v_1 = cp0_tlb_write_data_v_1; // @[myCPU.scala 974:32]
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 560:36]
      pre_decoder_branchD_flag <= 1'h0;
    end else if (_cfu_io_FlushD) begin // @[myCPU.scala 560:66]
      pre_decoder_branchD_flag <= 1'h0;
    end else if (_PCSrcD_T_1) begin
      pre_decoder_branchD_flag <= fifo_io_read_out_0[125];
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 562:34]
      pre_decoder_branchdata <= 6'h0;
    end else if (_pre_decoder_branchD_flag_T) begin // @[myCPU.scala 562:64]
      pre_decoder_branchdata <= 6'h0;
    end else if (_PCSrcD_T_1) begin
      pre_decoder_branchdata <= fifo_io_read_out_0[132:127];
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 561:28]
      pre_decoder_jump <= 1'h0;
    end else if (_pre_decoder_branchD_flag_T) begin // @[myCPU.scala 561:58]
      pre_decoder_jump <= 1'h0;
    end else if (_PCSrcD_T_1) begin
      pre_decoder_jump <= fifo_io_read_out_0[126];
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 563:26]
      pre_decoder_jr <= 1'h0;
    end else if (_pre_decoder_branchD_flag_T) begin // @[myCPU.scala 563:56]
      pre_decoder_jr <= 1'h0;
    end else if (_PCSrcD_T_1) begin
      pre_decoder_jr <= fifo_io_read_out_0[133];
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 931:25]
      resultE2M_Reg <= 32'h0;
    end else if (_mem_exception_T) begin // @[myCPU.scala 931:55]
      resultE2M_Reg <= 32'h0; // @[Mux.scala 101:{16,16} 81:58]
    end else if (_mem_exception_T_1) begin
      if (CP0ToRegE) begin
        if (2'h2 == _cfu_io_ForwardCP0E) begin
          resultE2M_Reg <= _mem2mem2_io_WriteCP0HiLoDataM;
        end else begin
          resultE2M_Reg <= _Forward_CP0_data_T_1;
        end
      end else if (_resultE_T_1) begin
        resultE2M_Reg <= _ex2mem_io_HiLoOutE;
      end else begin
        resultE2M_Reg <= _resultE_T_5;
      end
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 990:24]
      ResultM2_Reg <= 32'h0;
    end else if (_mem2_exception_T) begin // @[myCPU.scala 990:55]
      ResultM2_Reg <= 32'h0;
    end else if (_mem2_exception_T_1) begin
      ResultM2_Reg <= resultE2M_Reg;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 277:19]
      PCW_Reg <= 32'h0;
    end else if (_mem22wb_io_PCW != 32'h0) begin
      PCW_Reg <= _mem22wb_io_PCW;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 278:20]
      slot_Reg <= 1'h0;
    end else if (_PCW_Reg_T) begin
      slot_Reg <= _mem22wb_io_InDelaySlotW;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 279:29]
      branchjump_Jr_Reg <= 2'h0;
    end else if (_PCW_Reg_T) begin
      branchjump_Jr_Reg <= _mem22wb_io_BranchJump_JrW;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 283:25]
      reg_pc <= 32'h0; // @[myCPU.scala 283:25]
    end else begin
      reg_pc <= _mem22wb_io_PCW; // @[myCPU.scala 284:12]
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 603:20]
      wb_exception <= 1'h0;
    end else if (_cfu_io_FlushW) begin // @[myCPU.scala 603:50]
      wb_exception <= 1'h0;
    end else if (_cfu_io_StallW) begin
      wb_exception <= _mem22wb_io_ExceptionTypeM != 32'h0;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 327:24]
      pc_next_wait <= 32'h0; // @[Mux.scala 101:{16,16} myCPU.scala 181:24 731:26 398:31]
    end else if (ready_to_branch | stage_fec_2_branch_answer) begin
      if (fifo_io_point_write_en) begin
        if (pre_decoder_jump) begin
          if (pre_decoder_jr) begin
            pc_next_wait <= BranchRsD;
          end else begin
            pc_next_wait <= _PCJumpD_T_3;
          end
        end else if (_PCSrcD_T_3) begin
          pc_next_wait <= PCBranchD;
        end else begin
          pc_next_wait <= _if2id_io_PCPlus8D;
        end
      end else if (stage_fec_2_branch_answer) begin
        pc_next_wait <= stage_fec_2_pre_target_0;
      end else begin
        pc_next_wait <= _stage_fec_1_pc_next_T_1;
      end
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 382:22]
      commit_bru_reg <= 1'h1;
    end else if (_commit_cache_reg_T & commit_bru_reg) begin
      commit_bru_reg <= ~_cu_io1_commit_cache_ins;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 490:40]
      stage_fec_2_stall_reg <= 1'h0; // @[myCPU.scala 490:40]
    end else begin
      stage_fec_2_stall_reg <= stage2_stall; // @[myCPU.scala 491:27]
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 462:29]
      stage_fec_2_valid <= 1'h0; // @[myCPU.scala 462:51]
    end else if (stage2_stall) begin
      if (fifo_io_point_write_en) begin
        stage_fec_2_valid <= access_stage1_sram_valid;
      end else begin
        stage_fec_2_valid <= stage_fec_1_valid;
      end
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 332:102]
      pc_req_wait <= 1'h0; // @[myCPU.scala 333:21]
    end else begin
      pc_req_wait <= ~inst_sram_en & _pc_next_wait_T & _stage_fec_2_branch_answer_T_8 | _GEN_0;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 342:28]
      exception_Pc_reg <= 32'h0;
    end else if (_stage_fec_2_branch_answer_T_7) begin
      exception_Pc_reg <= _cp0_io_return_pc;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 347:58]
      returnPc_req_wait <= 1'h0; // @[myCPU.scala 348:27]
    end else begin
      returnPc_req_wait <= _T_4 & _stage_fec_2_branch_answer_T_7 | _GEN_2;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 381:24]
      commit_cache_reg <= 1'h1;
    end else if (_cfu_io_StallE & _cu_io1_commit_cache_ins) begin
      commit_cache_reg <= ~commit_cache_reg;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 444:29]
      stage_fec_1_valid <= 1'h0;
    end else begin
      stage_fec_1_valid <= stage2_stall | _stage_fec_1_valid_T_1;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 474:30]
      stage_fec_2_bht_0 <= 7'h0;
    end else if (stage2_flush) begin // @[myCPU.scala 474:51]
      stage_fec_2_bht_0 <= 7'h0;
    end else if (stage2_stall) begin
      stage_fec_2_bht_0 <= branch_prediction_with_blockram_io_bht_L;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 486:36]
      stage_fec_2_hascode_0 <= 4'h0;
    end else if (stage2_flush) begin // @[myCPU.scala 486:57]
      stage_fec_2_hascode_0 <= 4'h0;
    end else if (stage2_stall) begin
      stage_fec_2_hascode_0 <= _stage_fec_2_hascode_0_T_1;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 567:92]
      InDelaySlotF <= 1'h0; // @[myCPU.scala 568:22]
    end else begin
      InDelaySlotF <= (pre_decoder_branchD_flag | pre_decoder_jump) & ~_cfu_io_StallF | _GEN_6;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 591:20]
      id_exception <= 1'h0;
    end else if (_pre_decoder_branchD_flag_T) begin // @[myCPU.scala 591:50]
      id_exception <= 1'h0;
    end else if (_PCSrcD_T_1) begin
      id_exception <= fifo_io_read_out_0[1:0] != 2'h0 | fifo_io_read_out_0[135:134] != 2'h0;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 594:20]
      ex_exception <= 1'h0;
    end else if (_cfu_io_FlushE) begin // @[myCPU.scala 594:50]
      ex_exception <= 1'h0;
    end else if (_commit_cache_reg_T) begin
      ex_exception <= _id2ex_io_ExceptionTypeD != 32'h0;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 597:21]
      mem_exception <= 1'h0;
    end else if (_cfu_io_FlushM) begin // @[myCPU.scala 597:51]
      mem_exception <= 1'h0;
    end else if (_cfu_io_StallM) begin
      mem_exception <= _ex2mem_io_ExceptionTypeE != 32'h0;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 600:22]
      mem2_exception <= 1'h0;
    end else if (_cfu_io_FlushM2) begin // @[myCPU.scala 600:53]
      mem2_exception <= 1'h0;
    end else if (_cfu_io_StallM2) begin
      mem2_exception <= _mem2mem2_io_ExceptionTypeE != 32'h0;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 650:28]
      id_true_branch_state <= 1'h0;
    end else if (_pre_decoder_branchD_flag_T) begin // @[myCPU.scala 650:58]
      id_true_branch_state <= 1'h0;
    end else if (_PCSrcD_T_1) begin
      id_true_branch_state <= fifo_io_read_out_0[116];
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 680:27]
      inst_tlb_exceptionE <= 1'h0;
    end else if (_ex_exception_T) begin // @[myCPU.scala 680:57]
      inst_tlb_exceptionE <= 1'h0;
    end else if (_commit_cache_reg_T) begin
      inst_tlb_exceptionE <= _if2id_io_ExceptionTypeD_Out != 2'h0;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 711:30]
      true_branch_stateE <= 1'h0;
    end else if (_ex_exception_T) begin // @[myCPU.scala 711:61]
      true_branch_stateE <= 1'h0;
    end else if (_commit_cache_reg_T) begin
      true_branch_stateE <= _T_61;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 758:25]
      int_instanceE <= 6'h0;
    end else if (_ex_exception_T) begin // @[myCPU.scala 758:55]
      int_instanceE <= 6'h0;
    end else if (_commit_cache_reg_T) begin
      int_instanceE <= int_with_timer_int;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 759:25]
      int_instanceM <= 6'h0;
    end else if (_mem_exception_T) begin // @[myCPU.scala 759:55]
      int_instanceM <= 6'h0;
    end else if (_mem_exception_T_1) begin
      int_instanceM <= int_instanceE;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 760:26]
      int_instanceM2 <= 6'h0;
    end else if (_mem2_exception_T) begin // @[myCPU.scala 760:57]
      int_instanceM2 <= 6'h0;
    end else if (_mem2_exception_T_1) begin
      int_instanceM2 <= int_instanceM;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 761:25]
      int_instanceW <= 6'h0;
    end else if (_wb_exception_T) begin // @[myCPU.scala 761:55]
      int_instanceW <= 6'h0;
    end else if (_wb_exception_T_1) begin
      int_instanceW <= int_instanceM2;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 807:27]
      inst_tlb_exceptionM <= 1'h0;
    end else if (_mem_exception_T) begin // @[myCPU.scala 807:57]
      inst_tlb_exceptionM <= 1'h0;
    end else if (_mem_exception_T_1) begin
      inst_tlb_exceptionM <= inst_tlb_exceptionE;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 821:33]
      RD1ForWardE_r <= 32'h0; // @[myCPU.scala 811:34]
    end else if (!(_commit_cache_reg_T)) begin // @[myCPU.scala 825:88]
      if ((_cfu_io_ForwardAE[0] | _cfu_io_ForwardAE[1]) & ~Forward_Lock1E) begin // @[myCPU.scala 811:34]
        if (2'h3 == _cfu_io_ForwardAE) begin
          RD1ForWardE_r <= ResultM2_Reg;
        end else if (2'h2 == _cfu_io_ForwardAE) begin
          RD1ForWardE_r <= resultE2M_Reg;
        end else begin
          RD1ForWardE_r <= _RD1ForWardE_p_T_1;
        end
      end
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 821:33]
      RD2ForWardE_r <= 32'h0; // @[myCPU.scala 812:34]
    end else if (!(_commit_cache_reg_T)) begin // @[myCPU.scala 829:87]
      if ((_cfu_io_ForwardBE[0] | _cfu_io_ForwardBE[1]) & ~Forward_Lock2E) begin // @[myCPU.scala 812:34]
        if (2'h3 == _cfu_io_ForwardBE) begin
          RD2ForWardE_r <= ResultM2_Reg;
        end else if (2'h2 == _cfu_io_ForwardBE) begin
          RD2ForWardE_r <= resultE2M_Reg;
        end else begin
          RD2ForWardE_r <= _RD2ForWardE_p_T_1;
        end
      end
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 821:33]
      Forward_Lock1E <= 1'h0; // @[myCPU.scala 822:24]
    end else if (_commit_cache_reg_T) begin // @[myCPU.scala 825:88]
      Forward_Lock1E <= 1'h0; // @[myCPU.scala 826:28]
    end else if ((_cfu_io_ForwardAE[0] | _cfu_io_ForwardAE[1]) & ~Forward_Lock1E) begin // @[myCPU.scala 813:34]
      Forward_Lock1E <= ~(_ex2mem_io_MemToRegM | _mem2mem2_io_MemToRegM);
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 821:33]
      Forward_Lock2E <= 1'h0; // @[myCPU.scala 823:24]
    end else if (_commit_cache_reg_T) begin // @[myCPU.scala 829:87]
      Forward_Lock2E <= 1'h0; // @[myCPU.scala 830:28]
    end else if ((_cfu_io_ForwardBE[0] | _cfu_io_ForwardBE[1]) & ~Forward_Lock2E) begin // @[myCPU.scala 814:34]
      Forward_Lock2E <= _Forward_Lock1E_T_3;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 1043:33]
      tlb_exception_cp0_writeM2 <= 1'h0;
    end else if (_mem2_exception_T) begin // @[myCPU.scala 1043:64]
      tlb_exception_cp0_writeM2 <= 1'h0;
    end else if (_mem2_exception_T_1) begin
      tlb_exception_cp0_writeM2 <= __mem2mem2_io1_WriteCP0AddrE_T_1;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 1044:33]
      tlb_exception_co0_writeW <= 1'h0;
    end else if (_wb_exception_T) begin // @[myCPU.scala 1044:63]
      tlb_exception_co0_writeW <= 1'h0;
    end else if (_wb_exception_T_1) begin
      tlb_exception_co0_writeW <= tlb_exception_cp0_writeM2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pre_decoder_branchD_flag = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  pre_decoder_branchdata = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  pre_decoder_jump = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  pre_decoder_jr = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  resultE2M_Reg = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  ResultM2_Reg = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  PCW_Reg = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  slot_Reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  branchjump_Jr_Reg = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  reg_pc = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  wb_exception = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  pc_next_wait = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  commit_bru_reg = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  stage_fec_2_stall_reg = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  stage_fec_2_valid = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  pc_req_wait = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  exception_Pc_reg = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  returnPc_req_wait = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  commit_cache_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  stage_fec_1_valid = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  stage_fec_2_bht_0 = _RAND_20[6:0];
  _RAND_21 = {1{`RANDOM}};
  stage_fec_2_hascode_0 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  InDelaySlotF = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  id_exception = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  ex_exception = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  mem_exception = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  mem2_exception = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  id_true_branch_state = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  inst_tlb_exceptionE = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  true_branch_stateE = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  int_instanceE = _RAND_30[5:0];
  _RAND_31 = {1{`RANDOM}};
  int_instanceM = _RAND_31[5:0];
  _RAND_32 = {1{`RANDOM}};
  int_instanceM2 = _RAND_32[5:0];
  _RAND_33 = {1{`RANDOM}};
  int_instanceW = _RAND_33[5:0];
  _RAND_34 = {1{`RANDOM}};
  inst_tlb_exceptionM = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  RD1ForWardE_r = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  RD2ForWardE_r = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  Forward_Lock1E = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  Forward_Lock2E = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  tlb_exception_cp0_writeM2 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  tlb_exception_co0_writeW = _RAND_40[0:0];
`endif // RANDOMIZE_REG_INIT
  if (_T_2) begin
    pre_decoder_branchD_flag = 1'h0;
  end
  if (_T_2) begin
    pre_decoder_branchdata = 6'h0;
  end
  if (_T_2) begin
    pre_decoder_jump = 1'h0;
  end
  if (_T_2) begin
    pre_decoder_jr = 1'h0;
  end
  if (_T_2) begin
    resultE2M_Reg = 32'h0;
  end
  if (_T_2) begin
    ResultM2_Reg = 32'h0;
  end
  if (_T_2) begin
    PCW_Reg = 32'h0;
  end
  if (_T_2) begin
    slot_Reg = 1'h0;
  end
  if (_T_2) begin
    branchjump_Jr_Reg = 2'h0;
  end
  if (_T_2) begin
    reg_pc = 32'h0;
  end
  if (_T_2) begin
    wb_exception = 1'h0;
  end
  if (_T_2) begin
    pc_next_wait = 32'h0;
  end
  if (_T_2) begin
    commit_bru_reg = 1'h1;
  end
  if (_T_2) begin
    stage_fec_2_stall_reg = 1'h0;
  end
  if (_T_2) begin
    stage_fec_2_valid = 1'h0;
  end
  if (_T_2) begin
    pc_req_wait = 1'h0;
  end
  if (_T_2) begin
    exception_Pc_reg = 32'h0;
  end
  if (_T_2) begin
    returnPc_req_wait = 1'h0;
  end
  if (_T_2) begin
    commit_cache_reg = 1'h1;
  end
  if (_T_2) begin
    stage_fec_1_valid = 1'h0;
  end
  if (_T_2) begin
    stage_fec_2_bht_0 = 7'h0;
  end
  if (_T_2) begin
    stage_fec_2_hascode_0 = 4'h0;
  end
  if (_T_2) begin
    InDelaySlotF = 1'h0;
  end
  if (_T_2) begin
    id_exception = 1'h0;
  end
  if (_T_2) begin
    ex_exception = 1'h0;
  end
  if (_T_2) begin
    mem_exception = 1'h0;
  end
  if (_T_2) begin
    mem2_exception = 1'h0;
  end
  if (_T_2) begin
    id_true_branch_state = 1'h0;
  end
  if (_T_2) begin
    inst_tlb_exceptionE = 1'h0;
  end
  if (_T_2) begin
    true_branch_stateE = 1'h0;
  end
  if (_T_2) begin
    int_instanceE = 6'h0;
  end
  if (_T_2) begin
    int_instanceM = 6'h0;
  end
  if (_T_2) begin
    int_instanceM2 = 6'h0;
  end
  if (_T_2) begin
    int_instanceW = 6'h0;
  end
  if (_T_2) begin
    inst_tlb_exceptionM = 1'h0;
  end
  if (_T_2) begin
    RD1ForWardE_r = 32'h0;
  end
  if (_T_2) begin
    RD2ForWardE_r = 32'h0;
  end
  if (_T_2) begin
    Forward_Lock1E = 1'h0;
  end
  if (_T_2) begin
    Forward_Lock2E = 1'h0;
  end
  if (_T_2) begin
    tlb_exception_cp0_writeM2 = 1'h0;
  end
  if (_T_2) begin
    tlb_exception_co0_writeW = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module icache_tag(
  input         clock,
  input         reset,
  input         io_wen,
  input  [20:0] io_wdata,
  input  [31:0] io_addr,
  output        io_hit,
  output        io_valid,
  input  [7:0]  io_asid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
`endif // RANDOMIZE_REG_INIT
  reg [20:0] tag_regs_0; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_1; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_2; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_3; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_4; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_5; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_6; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_7; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_8; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_9; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_10; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_11; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_12; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_13; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_14; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_15; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_16; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_17; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_18; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_19; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_20; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_21; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_22; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_23; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_24; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_25; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_26; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_27; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_28; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_29; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_30; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_31; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_32; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_33; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_34; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_35; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_36; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_37; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_38; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_39; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_40; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_41; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_42; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_43; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_44; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_45; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_46; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_47; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_48; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_49; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_50; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_51; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_52; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_53; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_54; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_55; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_56; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_57; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_58; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_59; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_60; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_61; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_62; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_63; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_64; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_65; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_66; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_67; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_68; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_69; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_70; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_71; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_72; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_73; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_74; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_75; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_76; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_77; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_78; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_79; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_80; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_81; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_82; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_83; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_84; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_85; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_86; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_87; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_88; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_89; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_90; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_91; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_92; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_93; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_94; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_95; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_96; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_97; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_98; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_99; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_100; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_101; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_102; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_103; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_104; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_105; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_106; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_107; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_108; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_109; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_110; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_111; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_112; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_113; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_114; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_115; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_116; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_117; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_118; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_119; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_120; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_121; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_122; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_123; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_124; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_125; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_126; // @[icache_tag.scala 20:27]
  reg [20:0] tag_regs_127; // @[icache_tag.scala 20:27]
  reg [7:0] tag_asid_regs_0; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_1; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_2; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_3; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_4; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_5; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_6; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_7; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_8; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_9; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_10; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_11; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_12; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_13; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_14; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_15; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_16; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_17; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_18; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_19; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_20; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_21; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_22; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_23; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_24; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_25; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_26; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_27; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_28; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_29; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_30; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_31; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_32; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_33; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_34; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_35; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_36; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_37; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_38; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_39; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_40; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_41; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_42; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_43; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_44; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_45; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_46; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_47; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_48; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_49; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_50; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_51; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_52; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_53; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_54; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_55; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_56; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_57; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_58; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_59; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_60; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_61; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_62; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_63; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_64; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_65; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_66; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_67; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_68; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_69; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_70; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_71; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_72; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_73; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_74; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_75; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_76; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_77; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_78; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_79; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_80; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_81; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_82; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_83; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_84; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_85; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_86; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_87; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_88; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_89; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_90; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_91; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_92; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_93; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_94; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_95; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_96; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_97; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_98; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_99; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_100; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_101; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_102; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_103; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_104; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_105; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_106; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_107; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_108; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_109; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_110; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_111; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_112; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_113; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_114; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_115; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_116; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_117; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_118; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_119; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_120; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_121; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_122; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_123; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_124; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_125; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_126; // @[icache_tag.scala 21:32]
  reg [7:0] tag_asid_regs_127; // @[icache_tag.scala 21:32]
  wire [20:0] _GEN_1 = 7'h1 == io_addr[11:5] ? tag_regs_1 : tag_regs_0; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_2 = 7'h2 == io_addr[11:5] ? tag_regs_2 : _GEN_1; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_3 = 7'h3 == io_addr[11:5] ? tag_regs_3 : _GEN_2; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_4 = 7'h4 == io_addr[11:5] ? tag_regs_4 : _GEN_3; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_5 = 7'h5 == io_addr[11:5] ? tag_regs_5 : _GEN_4; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_6 = 7'h6 == io_addr[11:5] ? tag_regs_6 : _GEN_5; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_7 = 7'h7 == io_addr[11:5] ? tag_regs_7 : _GEN_6; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_8 = 7'h8 == io_addr[11:5] ? tag_regs_8 : _GEN_7; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_9 = 7'h9 == io_addr[11:5] ? tag_regs_9 : _GEN_8; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_10 = 7'ha == io_addr[11:5] ? tag_regs_10 : _GEN_9; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_11 = 7'hb == io_addr[11:5] ? tag_regs_11 : _GEN_10; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_12 = 7'hc == io_addr[11:5] ? tag_regs_12 : _GEN_11; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_13 = 7'hd == io_addr[11:5] ? tag_regs_13 : _GEN_12; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_14 = 7'he == io_addr[11:5] ? tag_regs_14 : _GEN_13; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_15 = 7'hf == io_addr[11:5] ? tag_regs_15 : _GEN_14; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_16 = 7'h10 == io_addr[11:5] ? tag_regs_16 : _GEN_15; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_17 = 7'h11 == io_addr[11:5] ? tag_regs_17 : _GEN_16; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_18 = 7'h12 == io_addr[11:5] ? tag_regs_18 : _GEN_17; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_19 = 7'h13 == io_addr[11:5] ? tag_regs_19 : _GEN_18; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_20 = 7'h14 == io_addr[11:5] ? tag_regs_20 : _GEN_19; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_21 = 7'h15 == io_addr[11:5] ? tag_regs_21 : _GEN_20; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_22 = 7'h16 == io_addr[11:5] ? tag_regs_22 : _GEN_21; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_23 = 7'h17 == io_addr[11:5] ? tag_regs_23 : _GEN_22; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_24 = 7'h18 == io_addr[11:5] ? tag_regs_24 : _GEN_23; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_25 = 7'h19 == io_addr[11:5] ? tag_regs_25 : _GEN_24; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_26 = 7'h1a == io_addr[11:5] ? tag_regs_26 : _GEN_25; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_27 = 7'h1b == io_addr[11:5] ? tag_regs_27 : _GEN_26; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_28 = 7'h1c == io_addr[11:5] ? tag_regs_28 : _GEN_27; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_29 = 7'h1d == io_addr[11:5] ? tag_regs_29 : _GEN_28; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_30 = 7'h1e == io_addr[11:5] ? tag_regs_30 : _GEN_29; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_31 = 7'h1f == io_addr[11:5] ? tag_regs_31 : _GEN_30; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_32 = 7'h20 == io_addr[11:5] ? tag_regs_32 : _GEN_31; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_33 = 7'h21 == io_addr[11:5] ? tag_regs_33 : _GEN_32; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_34 = 7'h22 == io_addr[11:5] ? tag_regs_34 : _GEN_33; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_35 = 7'h23 == io_addr[11:5] ? tag_regs_35 : _GEN_34; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_36 = 7'h24 == io_addr[11:5] ? tag_regs_36 : _GEN_35; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_37 = 7'h25 == io_addr[11:5] ? tag_regs_37 : _GEN_36; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_38 = 7'h26 == io_addr[11:5] ? tag_regs_38 : _GEN_37; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_39 = 7'h27 == io_addr[11:5] ? tag_regs_39 : _GEN_38; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_40 = 7'h28 == io_addr[11:5] ? tag_regs_40 : _GEN_39; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_41 = 7'h29 == io_addr[11:5] ? tag_regs_41 : _GEN_40; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_42 = 7'h2a == io_addr[11:5] ? tag_regs_42 : _GEN_41; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_43 = 7'h2b == io_addr[11:5] ? tag_regs_43 : _GEN_42; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_44 = 7'h2c == io_addr[11:5] ? tag_regs_44 : _GEN_43; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_45 = 7'h2d == io_addr[11:5] ? tag_regs_45 : _GEN_44; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_46 = 7'h2e == io_addr[11:5] ? tag_regs_46 : _GEN_45; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_47 = 7'h2f == io_addr[11:5] ? tag_regs_47 : _GEN_46; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_48 = 7'h30 == io_addr[11:5] ? tag_regs_48 : _GEN_47; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_49 = 7'h31 == io_addr[11:5] ? tag_regs_49 : _GEN_48; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_50 = 7'h32 == io_addr[11:5] ? tag_regs_50 : _GEN_49; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_51 = 7'h33 == io_addr[11:5] ? tag_regs_51 : _GEN_50; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_52 = 7'h34 == io_addr[11:5] ? tag_regs_52 : _GEN_51; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_53 = 7'h35 == io_addr[11:5] ? tag_regs_53 : _GEN_52; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_54 = 7'h36 == io_addr[11:5] ? tag_regs_54 : _GEN_53; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_55 = 7'h37 == io_addr[11:5] ? tag_regs_55 : _GEN_54; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_56 = 7'h38 == io_addr[11:5] ? tag_regs_56 : _GEN_55; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_57 = 7'h39 == io_addr[11:5] ? tag_regs_57 : _GEN_56; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_58 = 7'h3a == io_addr[11:5] ? tag_regs_58 : _GEN_57; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_59 = 7'h3b == io_addr[11:5] ? tag_regs_59 : _GEN_58; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_60 = 7'h3c == io_addr[11:5] ? tag_regs_60 : _GEN_59; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_61 = 7'h3d == io_addr[11:5] ? tag_regs_61 : _GEN_60; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_62 = 7'h3e == io_addr[11:5] ? tag_regs_62 : _GEN_61; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_63 = 7'h3f == io_addr[11:5] ? tag_regs_63 : _GEN_62; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_64 = 7'h40 == io_addr[11:5] ? tag_regs_64 : _GEN_63; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_65 = 7'h41 == io_addr[11:5] ? tag_regs_65 : _GEN_64; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_66 = 7'h42 == io_addr[11:5] ? tag_regs_66 : _GEN_65; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_67 = 7'h43 == io_addr[11:5] ? tag_regs_67 : _GEN_66; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_68 = 7'h44 == io_addr[11:5] ? tag_regs_68 : _GEN_67; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_69 = 7'h45 == io_addr[11:5] ? tag_regs_69 : _GEN_68; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_70 = 7'h46 == io_addr[11:5] ? tag_regs_70 : _GEN_69; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_71 = 7'h47 == io_addr[11:5] ? tag_regs_71 : _GEN_70; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_72 = 7'h48 == io_addr[11:5] ? tag_regs_72 : _GEN_71; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_73 = 7'h49 == io_addr[11:5] ? tag_regs_73 : _GEN_72; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_74 = 7'h4a == io_addr[11:5] ? tag_regs_74 : _GEN_73; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_75 = 7'h4b == io_addr[11:5] ? tag_regs_75 : _GEN_74; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_76 = 7'h4c == io_addr[11:5] ? tag_regs_76 : _GEN_75; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_77 = 7'h4d == io_addr[11:5] ? tag_regs_77 : _GEN_76; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_78 = 7'h4e == io_addr[11:5] ? tag_regs_78 : _GEN_77; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_79 = 7'h4f == io_addr[11:5] ? tag_regs_79 : _GEN_78; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_80 = 7'h50 == io_addr[11:5] ? tag_regs_80 : _GEN_79; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_81 = 7'h51 == io_addr[11:5] ? tag_regs_81 : _GEN_80; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_82 = 7'h52 == io_addr[11:5] ? tag_regs_82 : _GEN_81; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_83 = 7'h53 == io_addr[11:5] ? tag_regs_83 : _GEN_82; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_84 = 7'h54 == io_addr[11:5] ? tag_regs_84 : _GEN_83; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_85 = 7'h55 == io_addr[11:5] ? tag_regs_85 : _GEN_84; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_86 = 7'h56 == io_addr[11:5] ? tag_regs_86 : _GEN_85; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_87 = 7'h57 == io_addr[11:5] ? tag_regs_87 : _GEN_86; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_88 = 7'h58 == io_addr[11:5] ? tag_regs_88 : _GEN_87; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_89 = 7'h59 == io_addr[11:5] ? tag_regs_89 : _GEN_88; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_90 = 7'h5a == io_addr[11:5] ? tag_regs_90 : _GEN_89; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_91 = 7'h5b == io_addr[11:5] ? tag_regs_91 : _GEN_90; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_92 = 7'h5c == io_addr[11:5] ? tag_regs_92 : _GEN_91; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_93 = 7'h5d == io_addr[11:5] ? tag_regs_93 : _GEN_92; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_94 = 7'h5e == io_addr[11:5] ? tag_regs_94 : _GEN_93; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_95 = 7'h5f == io_addr[11:5] ? tag_regs_95 : _GEN_94; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_96 = 7'h60 == io_addr[11:5] ? tag_regs_96 : _GEN_95; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_97 = 7'h61 == io_addr[11:5] ? tag_regs_97 : _GEN_96; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_98 = 7'h62 == io_addr[11:5] ? tag_regs_98 : _GEN_97; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_99 = 7'h63 == io_addr[11:5] ? tag_regs_99 : _GEN_98; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_100 = 7'h64 == io_addr[11:5] ? tag_regs_100 : _GEN_99; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_101 = 7'h65 == io_addr[11:5] ? tag_regs_101 : _GEN_100; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_102 = 7'h66 == io_addr[11:5] ? tag_regs_102 : _GEN_101; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_103 = 7'h67 == io_addr[11:5] ? tag_regs_103 : _GEN_102; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_104 = 7'h68 == io_addr[11:5] ? tag_regs_104 : _GEN_103; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_105 = 7'h69 == io_addr[11:5] ? tag_regs_105 : _GEN_104; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_106 = 7'h6a == io_addr[11:5] ? tag_regs_106 : _GEN_105; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_107 = 7'h6b == io_addr[11:5] ? tag_regs_107 : _GEN_106; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_108 = 7'h6c == io_addr[11:5] ? tag_regs_108 : _GEN_107; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_109 = 7'h6d == io_addr[11:5] ? tag_regs_109 : _GEN_108; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_110 = 7'h6e == io_addr[11:5] ? tag_regs_110 : _GEN_109; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_111 = 7'h6f == io_addr[11:5] ? tag_regs_111 : _GEN_110; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_112 = 7'h70 == io_addr[11:5] ? tag_regs_112 : _GEN_111; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_113 = 7'h71 == io_addr[11:5] ? tag_regs_113 : _GEN_112; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_114 = 7'h72 == io_addr[11:5] ? tag_regs_114 : _GEN_113; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_115 = 7'h73 == io_addr[11:5] ? tag_regs_115 : _GEN_114; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_116 = 7'h74 == io_addr[11:5] ? tag_regs_116 : _GEN_115; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_117 = 7'h75 == io_addr[11:5] ? tag_regs_117 : _GEN_116; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_118 = 7'h76 == io_addr[11:5] ? tag_regs_118 : _GEN_117; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_119 = 7'h77 == io_addr[11:5] ? tag_regs_119 : _GEN_118; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_120 = 7'h78 == io_addr[11:5] ? tag_regs_120 : _GEN_119; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_121 = 7'h79 == io_addr[11:5] ? tag_regs_121 : _GEN_120; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_122 = 7'h7a == io_addr[11:5] ? tag_regs_122 : _GEN_121; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_123 = 7'h7b == io_addr[11:5] ? tag_regs_123 : _GEN_122; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_124 = 7'h7c == io_addr[11:5] ? tag_regs_124 : _GEN_123; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_125 = 7'h7d == io_addr[11:5] ? tag_regs_125 : _GEN_124; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_126 = 7'h7e == io_addr[11:5] ? tag_regs_126 : _GEN_125; // @[icache_tag.scala 24:{35,35}]
  wire [20:0] _GEN_127 = 7'h7f == io_addr[11:5] ? tag_regs_127 : _GEN_126; // @[icache_tag.scala 24:{35,35}]
  wire [7:0] _GEN_257 = 7'h1 == io_addr[11:5] ? tag_asid_regs_1 : tag_asid_regs_0; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_258 = 7'h2 == io_addr[11:5] ? tag_asid_regs_2 : _GEN_257; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_259 = 7'h3 == io_addr[11:5] ? tag_asid_regs_3 : _GEN_258; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_260 = 7'h4 == io_addr[11:5] ? tag_asid_regs_4 : _GEN_259; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_261 = 7'h5 == io_addr[11:5] ? tag_asid_regs_5 : _GEN_260; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_262 = 7'h6 == io_addr[11:5] ? tag_asid_regs_6 : _GEN_261; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_263 = 7'h7 == io_addr[11:5] ? tag_asid_regs_7 : _GEN_262; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_264 = 7'h8 == io_addr[11:5] ? tag_asid_regs_8 : _GEN_263; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_265 = 7'h9 == io_addr[11:5] ? tag_asid_regs_9 : _GEN_264; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_266 = 7'ha == io_addr[11:5] ? tag_asid_regs_10 : _GEN_265; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_267 = 7'hb == io_addr[11:5] ? tag_asid_regs_11 : _GEN_266; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_268 = 7'hc == io_addr[11:5] ? tag_asid_regs_12 : _GEN_267; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_269 = 7'hd == io_addr[11:5] ? tag_asid_regs_13 : _GEN_268; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_270 = 7'he == io_addr[11:5] ? tag_asid_regs_14 : _GEN_269; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_271 = 7'hf == io_addr[11:5] ? tag_asid_regs_15 : _GEN_270; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_272 = 7'h10 == io_addr[11:5] ? tag_asid_regs_16 : _GEN_271; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_273 = 7'h11 == io_addr[11:5] ? tag_asid_regs_17 : _GEN_272; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_274 = 7'h12 == io_addr[11:5] ? tag_asid_regs_18 : _GEN_273; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_275 = 7'h13 == io_addr[11:5] ? tag_asid_regs_19 : _GEN_274; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_276 = 7'h14 == io_addr[11:5] ? tag_asid_regs_20 : _GEN_275; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_277 = 7'h15 == io_addr[11:5] ? tag_asid_regs_21 : _GEN_276; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_278 = 7'h16 == io_addr[11:5] ? tag_asid_regs_22 : _GEN_277; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_279 = 7'h17 == io_addr[11:5] ? tag_asid_regs_23 : _GEN_278; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_280 = 7'h18 == io_addr[11:5] ? tag_asid_regs_24 : _GEN_279; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_281 = 7'h19 == io_addr[11:5] ? tag_asid_regs_25 : _GEN_280; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_282 = 7'h1a == io_addr[11:5] ? tag_asid_regs_26 : _GEN_281; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_283 = 7'h1b == io_addr[11:5] ? tag_asid_regs_27 : _GEN_282; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_284 = 7'h1c == io_addr[11:5] ? tag_asid_regs_28 : _GEN_283; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_285 = 7'h1d == io_addr[11:5] ? tag_asid_regs_29 : _GEN_284; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_286 = 7'h1e == io_addr[11:5] ? tag_asid_regs_30 : _GEN_285; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_287 = 7'h1f == io_addr[11:5] ? tag_asid_regs_31 : _GEN_286; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_288 = 7'h20 == io_addr[11:5] ? tag_asid_regs_32 : _GEN_287; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_289 = 7'h21 == io_addr[11:5] ? tag_asid_regs_33 : _GEN_288; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_290 = 7'h22 == io_addr[11:5] ? tag_asid_regs_34 : _GEN_289; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_291 = 7'h23 == io_addr[11:5] ? tag_asid_regs_35 : _GEN_290; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_292 = 7'h24 == io_addr[11:5] ? tag_asid_regs_36 : _GEN_291; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_293 = 7'h25 == io_addr[11:5] ? tag_asid_regs_37 : _GEN_292; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_294 = 7'h26 == io_addr[11:5] ? tag_asid_regs_38 : _GEN_293; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_295 = 7'h27 == io_addr[11:5] ? tag_asid_regs_39 : _GEN_294; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_296 = 7'h28 == io_addr[11:5] ? tag_asid_regs_40 : _GEN_295; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_297 = 7'h29 == io_addr[11:5] ? tag_asid_regs_41 : _GEN_296; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_298 = 7'h2a == io_addr[11:5] ? tag_asid_regs_42 : _GEN_297; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_299 = 7'h2b == io_addr[11:5] ? tag_asid_regs_43 : _GEN_298; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_300 = 7'h2c == io_addr[11:5] ? tag_asid_regs_44 : _GEN_299; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_301 = 7'h2d == io_addr[11:5] ? tag_asid_regs_45 : _GEN_300; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_302 = 7'h2e == io_addr[11:5] ? tag_asid_regs_46 : _GEN_301; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_303 = 7'h2f == io_addr[11:5] ? tag_asid_regs_47 : _GEN_302; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_304 = 7'h30 == io_addr[11:5] ? tag_asid_regs_48 : _GEN_303; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_305 = 7'h31 == io_addr[11:5] ? tag_asid_regs_49 : _GEN_304; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_306 = 7'h32 == io_addr[11:5] ? tag_asid_regs_50 : _GEN_305; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_307 = 7'h33 == io_addr[11:5] ? tag_asid_regs_51 : _GEN_306; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_308 = 7'h34 == io_addr[11:5] ? tag_asid_regs_52 : _GEN_307; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_309 = 7'h35 == io_addr[11:5] ? tag_asid_regs_53 : _GEN_308; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_310 = 7'h36 == io_addr[11:5] ? tag_asid_regs_54 : _GEN_309; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_311 = 7'h37 == io_addr[11:5] ? tag_asid_regs_55 : _GEN_310; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_312 = 7'h38 == io_addr[11:5] ? tag_asid_regs_56 : _GEN_311; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_313 = 7'h39 == io_addr[11:5] ? tag_asid_regs_57 : _GEN_312; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_314 = 7'h3a == io_addr[11:5] ? tag_asid_regs_58 : _GEN_313; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_315 = 7'h3b == io_addr[11:5] ? tag_asid_regs_59 : _GEN_314; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_316 = 7'h3c == io_addr[11:5] ? tag_asid_regs_60 : _GEN_315; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_317 = 7'h3d == io_addr[11:5] ? tag_asid_regs_61 : _GEN_316; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_318 = 7'h3e == io_addr[11:5] ? tag_asid_regs_62 : _GEN_317; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_319 = 7'h3f == io_addr[11:5] ? tag_asid_regs_63 : _GEN_318; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_320 = 7'h40 == io_addr[11:5] ? tag_asid_regs_64 : _GEN_319; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_321 = 7'h41 == io_addr[11:5] ? tag_asid_regs_65 : _GEN_320; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_322 = 7'h42 == io_addr[11:5] ? tag_asid_regs_66 : _GEN_321; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_323 = 7'h43 == io_addr[11:5] ? tag_asid_regs_67 : _GEN_322; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_324 = 7'h44 == io_addr[11:5] ? tag_asid_regs_68 : _GEN_323; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_325 = 7'h45 == io_addr[11:5] ? tag_asid_regs_69 : _GEN_324; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_326 = 7'h46 == io_addr[11:5] ? tag_asid_regs_70 : _GEN_325; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_327 = 7'h47 == io_addr[11:5] ? tag_asid_regs_71 : _GEN_326; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_328 = 7'h48 == io_addr[11:5] ? tag_asid_regs_72 : _GEN_327; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_329 = 7'h49 == io_addr[11:5] ? tag_asid_regs_73 : _GEN_328; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_330 = 7'h4a == io_addr[11:5] ? tag_asid_regs_74 : _GEN_329; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_331 = 7'h4b == io_addr[11:5] ? tag_asid_regs_75 : _GEN_330; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_332 = 7'h4c == io_addr[11:5] ? tag_asid_regs_76 : _GEN_331; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_333 = 7'h4d == io_addr[11:5] ? tag_asid_regs_77 : _GEN_332; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_334 = 7'h4e == io_addr[11:5] ? tag_asid_regs_78 : _GEN_333; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_335 = 7'h4f == io_addr[11:5] ? tag_asid_regs_79 : _GEN_334; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_336 = 7'h50 == io_addr[11:5] ? tag_asid_regs_80 : _GEN_335; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_337 = 7'h51 == io_addr[11:5] ? tag_asid_regs_81 : _GEN_336; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_338 = 7'h52 == io_addr[11:5] ? tag_asid_regs_82 : _GEN_337; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_339 = 7'h53 == io_addr[11:5] ? tag_asid_regs_83 : _GEN_338; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_340 = 7'h54 == io_addr[11:5] ? tag_asid_regs_84 : _GEN_339; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_341 = 7'h55 == io_addr[11:5] ? tag_asid_regs_85 : _GEN_340; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_342 = 7'h56 == io_addr[11:5] ? tag_asid_regs_86 : _GEN_341; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_343 = 7'h57 == io_addr[11:5] ? tag_asid_regs_87 : _GEN_342; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_344 = 7'h58 == io_addr[11:5] ? tag_asid_regs_88 : _GEN_343; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_345 = 7'h59 == io_addr[11:5] ? tag_asid_regs_89 : _GEN_344; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_346 = 7'h5a == io_addr[11:5] ? tag_asid_regs_90 : _GEN_345; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_347 = 7'h5b == io_addr[11:5] ? tag_asid_regs_91 : _GEN_346; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_348 = 7'h5c == io_addr[11:5] ? tag_asid_regs_92 : _GEN_347; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_349 = 7'h5d == io_addr[11:5] ? tag_asid_regs_93 : _GEN_348; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_350 = 7'h5e == io_addr[11:5] ? tag_asid_regs_94 : _GEN_349; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_351 = 7'h5f == io_addr[11:5] ? tag_asid_regs_95 : _GEN_350; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_352 = 7'h60 == io_addr[11:5] ? tag_asid_regs_96 : _GEN_351; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_353 = 7'h61 == io_addr[11:5] ? tag_asid_regs_97 : _GEN_352; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_354 = 7'h62 == io_addr[11:5] ? tag_asid_regs_98 : _GEN_353; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_355 = 7'h63 == io_addr[11:5] ? tag_asid_regs_99 : _GEN_354; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_356 = 7'h64 == io_addr[11:5] ? tag_asid_regs_100 : _GEN_355; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_357 = 7'h65 == io_addr[11:5] ? tag_asid_regs_101 : _GEN_356; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_358 = 7'h66 == io_addr[11:5] ? tag_asid_regs_102 : _GEN_357; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_359 = 7'h67 == io_addr[11:5] ? tag_asid_regs_103 : _GEN_358; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_360 = 7'h68 == io_addr[11:5] ? tag_asid_regs_104 : _GEN_359; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_361 = 7'h69 == io_addr[11:5] ? tag_asid_regs_105 : _GEN_360; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_362 = 7'h6a == io_addr[11:5] ? tag_asid_regs_106 : _GEN_361; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_363 = 7'h6b == io_addr[11:5] ? tag_asid_regs_107 : _GEN_362; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_364 = 7'h6c == io_addr[11:5] ? tag_asid_regs_108 : _GEN_363; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_365 = 7'h6d == io_addr[11:5] ? tag_asid_regs_109 : _GEN_364; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_366 = 7'h6e == io_addr[11:5] ? tag_asid_regs_110 : _GEN_365; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_367 = 7'h6f == io_addr[11:5] ? tag_asid_regs_111 : _GEN_366; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_368 = 7'h70 == io_addr[11:5] ? tag_asid_regs_112 : _GEN_367; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_369 = 7'h71 == io_addr[11:5] ? tag_asid_regs_113 : _GEN_368; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_370 = 7'h72 == io_addr[11:5] ? tag_asid_regs_114 : _GEN_369; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_371 = 7'h73 == io_addr[11:5] ? tag_asid_regs_115 : _GEN_370; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_372 = 7'h74 == io_addr[11:5] ? tag_asid_regs_116 : _GEN_371; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_373 = 7'h75 == io_addr[11:5] ? tag_asid_regs_117 : _GEN_372; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_374 = 7'h76 == io_addr[11:5] ? tag_asid_regs_118 : _GEN_373; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_375 = 7'h77 == io_addr[11:5] ? tag_asid_regs_119 : _GEN_374; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_376 = 7'h78 == io_addr[11:5] ? tag_asid_regs_120 : _GEN_375; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_377 = 7'h79 == io_addr[11:5] ? tag_asid_regs_121 : _GEN_376; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_378 = 7'h7a == io_addr[11:5] ? tag_asid_regs_122 : _GEN_377; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_379 = 7'h7b == io_addr[11:5] ? tag_asid_regs_123 : _GEN_378; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_380 = 7'h7c == io_addr[11:5] ? tag_asid_regs_124 : _GEN_379; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_381 = 7'h7d == io_addr[11:5] ? tag_asid_regs_125 : _GEN_380; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_382 = 7'h7e == io_addr[11:5] ? tag_asid_regs_126 : _GEN_381; // @[icache_tag.scala 25:{40,40}]
  wire [7:0] _GEN_383 = 7'h7f == io_addr[11:5] ? tag_asid_regs_127 : _GEN_382; // @[icache_tag.scala 25:{40,40}]
  assign io_hit = _GEN_127[19:0] == io_addr[31:12] & _GEN_383 == io_asid; // @[icache_tag.scala 29:50]
  assign io_valid = _GEN_127[20]; // @[icache_tag.scala 28:22]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_0 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h0 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_0 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_0 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_0 <= tag_regs_126;
      end else begin
        tag_regs_0 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_1 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h1 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_1 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_1 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_1 <= tag_regs_126;
      end else begin
        tag_regs_1 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_2 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h2 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_2 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_2 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_2 <= tag_regs_126;
      end else begin
        tag_regs_2 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_3 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h3 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_3 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_3 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_3 <= tag_regs_126;
      end else begin
        tag_regs_3 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_4 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h4 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_4 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_4 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_4 <= tag_regs_126;
      end else begin
        tag_regs_4 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_5 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h5 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_5 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_5 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_5 <= tag_regs_126;
      end else begin
        tag_regs_5 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_6 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h6 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_6 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_6 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_6 <= tag_regs_126;
      end else begin
        tag_regs_6 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_7 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h7 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_7 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_7 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_7 <= tag_regs_126;
      end else begin
        tag_regs_7 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_8 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h8 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_8 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_8 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_8 <= tag_regs_126;
      end else begin
        tag_regs_8 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_9 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h9 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_9 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_9 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_9 <= tag_regs_126;
      end else begin
        tag_regs_9 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_10 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'ha == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_10 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_10 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_10 <= tag_regs_126;
      end else begin
        tag_regs_10 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_11 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'hb == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_11 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_11 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_11 <= tag_regs_126;
      end else begin
        tag_regs_11 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_12 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'hc == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_12 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_12 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_12 <= tag_regs_126;
      end else begin
        tag_regs_12 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_13 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'hd == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_13 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_13 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_13 <= tag_regs_126;
      end else begin
        tag_regs_13 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_14 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'he == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_14 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_14 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_14 <= tag_regs_126;
      end else begin
        tag_regs_14 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_15 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'hf == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_15 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_15 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_15 <= tag_regs_126;
      end else begin
        tag_regs_15 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_16 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h10 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_16 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_16 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_16 <= tag_regs_126;
      end else begin
        tag_regs_16 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_17 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h11 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_17 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_17 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_17 <= tag_regs_126;
      end else begin
        tag_regs_17 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_18 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h12 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_18 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_18 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_18 <= tag_regs_126;
      end else begin
        tag_regs_18 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_19 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h13 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_19 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_19 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_19 <= tag_regs_126;
      end else begin
        tag_regs_19 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_20 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h14 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_20 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_20 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_20 <= tag_regs_126;
      end else begin
        tag_regs_20 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_21 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h15 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_21 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_21 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_21 <= tag_regs_126;
      end else begin
        tag_regs_21 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_22 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h16 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_22 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_22 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_22 <= tag_regs_126;
      end else begin
        tag_regs_22 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_23 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h17 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_23 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_23 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_23 <= tag_regs_126;
      end else begin
        tag_regs_23 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_24 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h18 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_24 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_24 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_24 <= tag_regs_126;
      end else begin
        tag_regs_24 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_25 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h19 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_25 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_25 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_25 <= tag_regs_126;
      end else begin
        tag_regs_25 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_26 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h1a == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_26 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_26 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_26 <= tag_regs_126;
      end else begin
        tag_regs_26 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_27 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h1b == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_27 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_27 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_27 <= tag_regs_126;
      end else begin
        tag_regs_27 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_28 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h1c == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_28 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_28 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_28 <= tag_regs_126;
      end else begin
        tag_regs_28 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_29 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h1d == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_29 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_29 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_29 <= tag_regs_126;
      end else begin
        tag_regs_29 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_30 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h1e == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_30 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_30 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_30 <= tag_regs_126;
      end else begin
        tag_regs_30 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_31 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h1f == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_31 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_31 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_31 <= tag_regs_126;
      end else begin
        tag_regs_31 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_32 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h20 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_32 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_32 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_32 <= tag_regs_126;
      end else begin
        tag_regs_32 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_33 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h21 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_33 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_33 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_33 <= tag_regs_126;
      end else begin
        tag_regs_33 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_34 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h22 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_34 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_34 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_34 <= tag_regs_126;
      end else begin
        tag_regs_34 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_35 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h23 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_35 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_35 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_35 <= tag_regs_126;
      end else begin
        tag_regs_35 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_36 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h24 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_36 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_36 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_36 <= tag_regs_126;
      end else begin
        tag_regs_36 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_37 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h25 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_37 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_37 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_37 <= tag_regs_126;
      end else begin
        tag_regs_37 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_38 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h26 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_38 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_38 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_38 <= tag_regs_126;
      end else begin
        tag_regs_38 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_39 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h27 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_39 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_39 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_39 <= tag_regs_126;
      end else begin
        tag_regs_39 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_40 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h28 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_40 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_40 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_40 <= tag_regs_126;
      end else begin
        tag_regs_40 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_41 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h29 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_41 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_41 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_41 <= tag_regs_126;
      end else begin
        tag_regs_41 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_42 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h2a == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_42 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_42 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_42 <= tag_regs_126;
      end else begin
        tag_regs_42 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_43 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h2b == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_43 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_43 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_43 <= tag_regs_126;
      end else begin
        tag_regs_43 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_44 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h2c == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_44 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_44 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_44 <= tag_regs_126;
      end else begin
        tag_regs_44 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_45 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h2d == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_45 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_45 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_45 <= tag_regs_126;
      end else begin
        tag_regs_45 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_46 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h2e == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_46 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_46 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_46 <= tag_regs_126;
      end else begin
        tag_regs_46 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_47 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h2f == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_47 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_47 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_47 <= tag_regs_126;
      end else begin
        tag_regs_47 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_48 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h30 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_48 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_48 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_48 <= tag_regs_126;
      end else begin
        tag_regs_48 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_49 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h31 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_49 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_49 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_49 <= tag_regs_126;
      end else begin
        tag_regs_49 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_50 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h32 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_50 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_50 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_50 <= tag_regs_126;
      end else begin
        tag_regs_50 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_51 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h33 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_51 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_51 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_51 <= tag_regs_126;
      end else begin
        tag_regs_51 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_52 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h34 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_52 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_52 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_52 <= tag_regs_126;
      end else begin
        tag_regs_52 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_53 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h35 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_53 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_53 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_53 <= tag_regs_126;
      end else begin
        tag_regs_53 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_54 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h36 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_54 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_54 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_54 <= tag_regs_126;
      end else begin
        tag_regs_54 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_55 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h37 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_55 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_55 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_55 <= tag_regs_126;
      end else begin
        tag_regs_55 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_56 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h38 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_56 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_56 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_56 <= tag_regs_126;
      end else begin
        tag_regs_56 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_57 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h39 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_57 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_57 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_57 <= tag_regs_126;
      end else begin
        tag_regs_57 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_58 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h3a == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_58 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_58 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_58 <= tag_regs_126;
      end else begin
        tag_regs_58 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_59 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h3b == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_59 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_59 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_59 <= tag_regs_126;
      end else begin
        tag_regs_59 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_60 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h3c == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_60 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_60 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_60 <= tag_regs_126;
      end else begin
        tag_regs_60 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_61 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h3d == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_61 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_61 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_61 <= tag_regs_126;
      end else begin
        tag_regs_61 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_62 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h3e == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_62 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_62 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_62 <= tag_regs_126;
      end else begin
        tag_regs_62 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_63 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h3f == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_63 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_63 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_63 <= tag_regs_126;
      end else begin
        tag_regs_63 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_64 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h40 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_64 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_64 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_64 <= tag_regs_126;
      end else begin
        tag_regs_64 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_65 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h41 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_65 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_65 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_65 <= tag_regs_126;
      end else begin
        tag_regs_65 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_66 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h42 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_66 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_66 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_66 <= tag_regs_126;
      end else begin
        tag_regs_66 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_67 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h43 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_67 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_67 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_67 <= tag_regs_126;
      end else begin
        tag_regs_67 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_68 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h44 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_68 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_68 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_68 <= tag_regs_126;
      end else begin
        tag_regs_68 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_69 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h45 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_69 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_69 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_69 <= tag_regs_126;
      end else begin
        tag_regs_69 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_70 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h46 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_70 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_70 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_70 <= tag_regs_126;
      end else begin
        tag_regs_70 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_71 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h47 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_71 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_71 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_71 <= tag_regs_126;
      end else begin
        tag_regs_71 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_72 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h48 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_72 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_72 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_72 <= tag_regs_126;
      end else begin
        tag_regs_72 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_73 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h49 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_73 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_73 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_73 <= tag_regs_126;
      end else begin
        tag_regs_73 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_74 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h4a == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_74 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_74 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_74 <= tag_regs_126;
      end else begin
        tag_regs_74 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_75 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h4b == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_75 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_75 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_75 <= tag_regs_126;
      end else begin
        tag_regs_75 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_76 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h4c == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_76 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_76 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_76 <= tag_regs_126;
      end else begin
        tag_regs_76 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_77 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h4d == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_77 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_77 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_77 <= tag_regs_126;
      end else begin
        tag_regs_77 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_78 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h4e == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_78 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_78 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_78 <= tag_regs_126;
      end else begin
        tag_regs_78 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_79 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h4f == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_79 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_79 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_79 <= tag_regs_126;
      end else begin
        tag_regs_79 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_80 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h50 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_80 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_80 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_80 <= tag_regs_126;
      end else begin
        tag_regs_80 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_81 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h51 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_81 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_81 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_81 <= tag_regs_126;
      end else begin
        tag_regs_81 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_82 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h52 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_82 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_82 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_82 <= tag_regs_126;
      end else begin
        tag_regs_82 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_83 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h53 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_83 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_83 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_83 <= tag_regs_126;
      end else begin
        tag_regs_83 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_84 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h54 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_84 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_84 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_84 <= tag_regs_126;
      end else begin
        tag_regs_84 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_85 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h55 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_85 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_85 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_85 <= tag_regs_126;
      end else begin
        tag_regs_85 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_86 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h56 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_86 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_86 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_86 <= tag_regs_126;
      end else begin
        tag_regs_86 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_87 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h57 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_87 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_87 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_87 <= tag_regs_126;
      end else begin
        tag_regs_87 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_88 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h58 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_88 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_88 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_88 <= tag_regs_126;
      end else begin
        tag_regs_88 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_89 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h59 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_89 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_89 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_89 <= tag_regs_126;
      end else begin
        tag_regs_89 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_90 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h5a == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_90 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_90 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_90 <= tag_regs_126;
      end else begin
        tag_regs_90 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_91 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h5b == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_91 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_91 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_91 <= tag_regs_126;
      end else begin
        tag_regs_91 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_92 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h5c == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_92 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_92 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_92 <= tag_regs_126;
      end else begin
        tag_regs_92 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_93 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h5d == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_93 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_93 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_93 <= tag_regs_126;
      end else begin
        tag_regs_93 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_94 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h5e == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_94 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_94 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_94 <= tag_regs_126;
      end else begin
        tag_regs_94 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_95 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h5f == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_95 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_95 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_95 <= tag_regs_126;
      end else begin
        tag_regs_95 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_96 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h60 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_96 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_96 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_96 <= tag_regs_126;
      end else begin
        tag_regs_96 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_97 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h61 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_97 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_97 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_97 <= tag_regs_126;
      end else begin
        tag_regs_97 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_98 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h62 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_98 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_98 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_98 <= tag_regs_126;
      end else begin
        tag_regs_98 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_99 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h63 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_99 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_99 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_99 <= tag_regs_126;
      end else begin
        tag_regs_99 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_100 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h64 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_100 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_100 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_100 <= tag_regs_126;
      end else begin
        tag_regs_100 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_101 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h65 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_101 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_101 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_101 <= tag_regs_126;
      end else begin
        tag_regs_101 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_102 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h66 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_102 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_102 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_102 <= tag_regs_126;
      end else begin
        tag_regs_102 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_103 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h67 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_103 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_103 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_103 <= tag_regs_126;
      end else begin
        tag_regs_103 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_104 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h68 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_104 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_104 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_104 <= tag_regs_126;
      end else begin
        tag_regs_104 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_105 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h69 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_105 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_105 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_105 <= tag_regs_126;
      end else begin
        tag_regs_105 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_106 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h6a == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_106 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_106 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_106 <= tag_regs_126;
      end else begin
        tag_regs_106 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_107 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h6b == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_107 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_107 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_107 <= tag_regs_126;
      end else begin
        tag_regs_107 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_108 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h6c == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_108 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_108 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_108 <= tag_regs_126;
      end else begin
        tag_regs_108 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_109 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h6d == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_109 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_109 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_109 <= tag_regs_126;
      end else begin
        tag_regs_109 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_110 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h6e == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_110 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_110 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_110 <= tag_regs_126;
      end else begin
        tag_regs_110 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_111 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h6f == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_111 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_111 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_111 <= tag_regs_126;
      end else begin
        tag_regs_111 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_112 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h70 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_112 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_112 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_112 <= tag_regs_126;
      end else begin
        tag_regs_112 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_113 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h71 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_113 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_113 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_113 <= tag_regs_126;
      end else begin
        tag_regs_113 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_114 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h72 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_114 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_114 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_114 <= tag_regs_126;
      end else begin
        tag_regs_114 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_115 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h73 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_115 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_115 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_115 <= tag_regs_126;
      end else begin
        tag_regs_115 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_116 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h74 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_116 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_116 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_116 <= tag_regs_126;
      end else begin
        tag_regs_116 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_117 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h75 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_117 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_117 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_117 <= tag_regs_126;
      end else begin
        tag_regs_117 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_118 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h76 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_118 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_118 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_118 <= tag_regs_126;
      end else begin
        tag_regs_118 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_119 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h77 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_119 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_119 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_119 <= tag_regs_126;
      end else begin
        tag_regs_119 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_120 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h78 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_120 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_120 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_120 <= tag_regs_126;
      end else begin
        tag_regs_120 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_121 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h79 == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_121 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_121 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_121 <= tag_regs_126;
      end else begin
        tag_regs_121 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_122 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h7a == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_122 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_122 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_122 <= tag_regs_126;
      end else begin
        tag_regs_122 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_123 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h7b == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_123 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_123 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_123 <= tag_regs_126;
      end else begin
        tag_regs_123 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_124 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h7c == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_124 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_124 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_124 <= tag_regs_126;
      end else begin
        tag_regs_124 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_125 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h7d == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_125 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_125 <= tag_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_regs_125 <= tag_regs_126;
      end else begin
        tag_regs_125 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_126 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h7e == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_126 <= io_wdata;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_regs_126 <= tag_regs_127;
      end else if (!(7'h7e == io_addr[11:5])) begin
        tag_regs_126 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 24:29]
      tag_regs_127 <= 21'h0; // @[icache_tag.scala 24:{35,35,35,35,35}]
    end else if (7'h7f == io_addr[11:5]) begin // @[icache_tag.scala 20:27]
      if (io_wen) begin
        tag_regs_127 <= io_wdata;
      end else if (!(7'h7f == io_addr[11:5])) begin
        if (7'h7e == io_addr[11:5]) begin
          tag_regs_127 <= tag_regs_126;
        end else begin
          tag_regs_127 <= _GEN_125;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_0 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h0 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_0 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_0 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_0 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_0 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_1 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h1 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_1 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_1 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_1 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_1 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_2 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h2 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_2 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_2 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_2 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_2 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_3 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h3 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_3 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_3 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_3 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_3 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_4 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h4 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_4 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_4 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_4 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_4 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_5 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h5 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_5 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_5 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_5 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_5 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_6 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h6 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_6 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_6 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_6 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_6 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_7 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h7 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_7 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_7 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_7 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_7 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_8 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h8 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_8 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_8 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_8 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_8 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_9 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h9 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_9 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_9 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_9 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_9 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_10 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'ha == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_10 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_10 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_10 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_10 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_11 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'hb == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_11 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_11 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_11 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_11 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_12 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'hc == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_12 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_12 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_12 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_12 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_13 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'hd == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_13 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_13 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_13 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_13 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_14 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'he == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_14 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_14 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_14 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_14 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_15 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'hf == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_15 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_15 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_15 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_15 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_16 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h10 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_16 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_16 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_16 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_16 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_17 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h11 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_17 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_17 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_17 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_17 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_18 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h12 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_18 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_18 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_18 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_18 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_19 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h13 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_19 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_19 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_19 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_19 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_20 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h14 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_20 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_20 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_20 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_20 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_21 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h15 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_21 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_21 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_21 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_21 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_22 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h16 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_22 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_22 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_22 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_22 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_23 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h17 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_23 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_23 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_23 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_23 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_24 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h18 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_24 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_24 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_24 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_24 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_25 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h19 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_25 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_25 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_25 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_25 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_26 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h1a == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_26 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_26 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_26 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_26 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_27 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h1b == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_27 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_27 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_27 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_27 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_28 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h1c == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_28 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_28 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_28 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_28 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_29 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h1d == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_29 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_29 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_29 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_29 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_30 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h1e == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_30 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_30 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_30 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_30 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_31 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h1f == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_31 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_31 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_31 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_31 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_32 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h20 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_32 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_32 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_32 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_32 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_33 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h21 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_33 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_33 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_33 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_33 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_34 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h22 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_34 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_34 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_34 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_34 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_35 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h23 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_35 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_35 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_35 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_35 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_36 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h24 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_36 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_36 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_36 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_36 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_37 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h25 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_37 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_37 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_37 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_37 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_38 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h26 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_38 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_38 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_38 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_38 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_39 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h27 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_39 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_39 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_39 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_39 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_40 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h28 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_40 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_40 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_40 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_40 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_41 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h29 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_41 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_41 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_41 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_41 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_42 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h2a == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_42 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_42 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_42 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_42 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_43 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h2b == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_43 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_43 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_43 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_43 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_44 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h2c == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_44 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_44 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_44 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_44 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_45 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h2d == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_45 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_45 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_45 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_45 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_46 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h2e == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_46 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_46 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_46 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_46 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_47 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h2f == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_47 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_47 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_47 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_47 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_48 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h30 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_48 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_48 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_48 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_48 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_49 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h31 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_49 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_49 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_49 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_49 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_50 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h32 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_50 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_50 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_50 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_50 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_51 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h33 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_51 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_51 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_51 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_51 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_52 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h34 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_52 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_52 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_52 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_52 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_53 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h35 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_53 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_53 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_53 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_53 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_54 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h36 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_54 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_54 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_54 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_54 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_55 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h37 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_55 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_55 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_55 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_55 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_56 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h38 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_56 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_56 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_56 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_56 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_57 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h39 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_57 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_57 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_57 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_57 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_58 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h3a == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_58 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_58 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_58 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_58 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_59 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h3b == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_59 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_59 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_59 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_59 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_60 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h3c == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_60 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_60 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_60 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_60 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_61 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h3d == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_61 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_61 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_61 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_61 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_62 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h3e == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_62 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_62 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_62 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_62 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_63 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h3f == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_63 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_63 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_63 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_63 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_64 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h40 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_64 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_64 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_64 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_64 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_65 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h41 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_65 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_65 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_65 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_65 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_66 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h42 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_66 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_66 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_66 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_66 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_67 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h43 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_67 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_67 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_67 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_67 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_68 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h44 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_68 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_68 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_68 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_68 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_69 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h45 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_69 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_69 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_69 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_69 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_70 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h46 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_70 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_70 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_70 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_70 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_71 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h47 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_71 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_71 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_71 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_71 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_72 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h48 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_72 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_72 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_72 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_72 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_73 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h49 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_73 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_73 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_73 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_73 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_74 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h4a == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_74 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_74 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_74 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_74 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_75 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h4b == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_75 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_75 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_75 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_75 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_76 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h4c == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_76 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_76 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_76 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_76 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_77 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h4d == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_77 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_77 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_77 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_77 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_78 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h4e == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_78 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_78 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_78 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_78 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_79 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h4f == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_79 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_79 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_79 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_79 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_80 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h50 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_80 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_80 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_80 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_80 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_81 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h51 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_81 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_81 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_81 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_81 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_82 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h52 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_82 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_82 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_82 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_82 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_83 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h53 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_83 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_83 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_83 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_83 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_84 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h54 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_84 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_84 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_84 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_84 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_85 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h55 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_85 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_85 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_85 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_85 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_86 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h56 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_86 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_86 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_86 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_86 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_87 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h57 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_87 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_87 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_87 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_87 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_88 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h58 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_88 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_88 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_88 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_88 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_89 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h59 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_89 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_89 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_89 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_89 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_90 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h5a == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_90 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_90 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_90 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_90 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_91 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h5b == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_91 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_91 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_91 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_91 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_92 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h5c == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_92 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_92 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_92 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_92 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_93 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h5d == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_93 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_93 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_93 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_93 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_94 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h5e == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_94 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_94 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_94 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_94 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_95 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h5f == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_95 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_95 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_95 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_95 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_96 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h60 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_96 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_96 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_96 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_96 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_97 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h61 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_97 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_97 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_97 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_97 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_98 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h62 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_98 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_98 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_98 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_98 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_99 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h63 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_99 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_99 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_99 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_99 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_100 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h64 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_100 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_100 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_100 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_100 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_101 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h65 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_101 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_101 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_101 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_101 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_102 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h66 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_102 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_102 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_102 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_102 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_103 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h67 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_103 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_103 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_103 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_103 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_104 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h68 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_104 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_104 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_104 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_104 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_105 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h69 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_105 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_105 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_105 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_105 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_106 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h6a == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_106 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_106 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_106 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_106 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_107 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h6b == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_107 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_107 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_107 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_107 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_108 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h6c == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_108 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_108 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_108 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_108 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_109 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h6d == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_109 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_109 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_109 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_109 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_110 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h6e == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_110 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_110 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_110 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_110 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_111 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h6f == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_111 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_111 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_111 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_111 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_112 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h70 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_112 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_112 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_112 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_112 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_113 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h71 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_113 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_113 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_113 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_113 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_114 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h72 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_114 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_114 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_114 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_114 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_115 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h73 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_115 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_115 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_115 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_115 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_116 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h74 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_116 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_116 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_116 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_116 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_117 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h75 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_117 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_117 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_117 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_117 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_118 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h76 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_118 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_118 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_118 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_118 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_119 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h77 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_119 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_119 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_119 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_119 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_120 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h78 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_120 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_120 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_120 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_120 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_121 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h79 == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_121 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_121 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_121 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_121 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_122 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h7a == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_122 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_122 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_122 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_122 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_123 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h7b == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_123 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_123 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_123 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_123 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_124 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h7c == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_124 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_124 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_124 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_124 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_125 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h7d == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_125 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_125 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[11:5]) begin
        tag_asid_regs_125 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_125 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_126 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h7e == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_126 <= io_asid;
      end else if (7'h7f == io_addr[11:5]) begin
        tag_asid_regs_126 <= tag_asid_regs_127;
      end else if (!(7'h7e == io_addr[11:5])) begin
        tag_asid_regs_126 <= _GEN_381;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 25:34]
      tag_asid_regs_127 <= 8'h0; // @[icache_tag.scala 25:{40,40,40,40,40}]
    end else if (7'h7f == io_addr[11:5]) begin // @[icache_tag.scala 21:32]
      if (io_wen) begin
        tag_asid_regs_127 <= io_asid;
      end else if (!(7'h7f == io_addr[11:5])) begin
        if (7'h7e == io_addr[11:5]) begin
          tag_asid_regs_127 <= tag_asid_regs_126;
        end else begin
          tag_asid_regs_127 <= _GEN_381;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_regs_0 = _RAND_0[20:0];
  _RAND_1 = {1{`RANDOM}};
  tag_regs_1 = _RAND_1[20:0];
  _RAND_2 = {1{`RANDOM}};
  tag_regs_2 = _RAND_2[20:0];
  _RAND_3 = {1{`RANDOM}};
  tag_regs_3 = _RAND_3[20:0];
  _RAND_4 = {1{`RANDOM}};
  tag_regs_4 = _RAND_4[20:0];
  _RAND_5 = {1{`RANDOM}};
  tag_regs_5 = _RAND_5[20:0];
  _RAND_6 = {1{`RANDOM}};
  tag_regs_6 = _RAND_6[20:0];
  _RAND_7 = {1{`RANDOM}};
  tag_regs_7 = _RAND_7[20:0];
  _RAND_8 = {1{`RANDOM}};
  tag_regs_8 = _RAND_8[20:0];
  _RAND_9 = {1{`RANDOM}};
  tag_regs_9 = _RAND_9[20:0];
  _RAND_10 = {1{`RANDOM}};
  tag_regs_10 = _RAND_10[20:0];
  _RAND_11 = {1{`RANDOM}};
  tag_regs_11 = _RAND_11[20:0];
  _RAND_12 = {1{`RANDOM}};
  tag_regs_12 = _RAND_12[20:0];
  _RAND_13 = {1{`RANDOM}};
  tag_regs_13 = _RAND_13[20:0];
  _RAND_14 = {1{`RANDOM}};
  tag_regs_14 = _RAND_14[20:0];
  _RAND_15 = {1{`RANDOM}};
  tag_regs_15 = _RAND_15[20:0];
  _RAND_16 = {1{`RANDOM}};
  tag_regs_16 = _RAND_16[20:0];
  _RAND_17 = {1{`RANDOM}};
  tag_regs_17 = _RAND_17[20:0];
  _RAND_18 = {1{`RANDOM}};
  tag_regs_18 = _RAND_18[20:0];
  _RAND_19 = {1{`RANDOM}};
  tag_regs_19 = _RAND_19[20:0];
  _RAND_20 = {1{`RANDOM}};
  tag_regs_20 = _RAND_20[20:0];
  _RAND_21 = {1{`RANDOM}};
  tag_regs_21 = _RAND_21[20:0];
  _RAND_22 = {1{`RANDOM}};
  tag_regs_22 = _RAND_22[20:0];
  _RAND_23 = {1{`RANDOM}};
  tag_regs_23 = _RAND_23[20:0];
  _RAND_24 = {1{`RANDOM}};
  tag_regs_24 = _RAND_24[20:0];
  _RAND_25 = {1{`RANDOM}};
  tag_regs_25 = _RAND_25[20:0];
  _RAND_26 = {1{`RANDOM}};
  tag_regs_26 = _RAND_26[20:0];
  _RAND_27 = {1{`RANDOM}};
  tag_regs_27 = _RAND_27[20:0];
  _RAND_28 = {1{`RANDOM}};
  tag_regs_28 = _RAND_28[20:0];
  _RAND_29 = {1{`RANDOM}};
  tag_regs_29 = _RAND_29[20:0];
  _RAND_30 = {1{`RANDOM}};
  tag_regs_30 = _RAND_30[20:0];
  _RAND_31 = {1{`RANDOM}};
  tag_regs_31 = _RAND_31[20:0];
  _RAND_32 = {1{`RANDOM}};
  tag_regs_32 = _RAND_32[20:0];
  _RAND_33 = {1{`RANDOM}};
  tag_regs_33 = _RAND_33[20:0];
  _RAND_34 = {1{`RANDOM}};
  tag_regs_34 = _RAND_34[20:0];
  _RAND_35 = {1{`RANDOM}};
  tag_regs_35 = _RAND_35[20:0];
  _RAND_36 = {1{`RANDOM}};
  tag_regs_36 = _RAND_36[20:0];
  _RAND_37 = {1{`RANDOM}};
  tag_regs_37 = _RAND_37[20:0];
  _RAND_38 = {1{`RANDOM}};
  tag_regs_38 = _RAND_38[20:0];
  _RAND_39 = {1{`RANDOM}};
  tag_regs_39 = _RAND_39[20:0];
  _RAND_40 = {1{`RANDOM}};
  tag_regs_40 = _RAND_40[20:0];
  _RAND_41 = {1{`RANDOM}};
  tag_regs_41 = _RAND_41[20:0];
  _RAND_42 = {1{`RANDOM}};
  tag_regs_42 = _RAND_42[20:0];
  _RAND_43 = {1{`RANDOM}};
  tag_regs_43 = _RAND_43[20:0];
  _RAND_44 = {1{`RANDOM}};
  tag_regs_44 = _RAND_44[20:0];
  _RAND_45 = {1{`RANDOM}};
  tag_regs_45 = _RAND_45[20:0];
  _RAND_46 = {1{`RANDOM}};
  tag_regs_46 = _RAND_46[20:0];
  _RAND_47 = {1{`RANDOM}};
  tag_regs_47 = _RAND_47[20:0];
  _RAND_48 = {1{`RANDOM}};
  tag_regs_48 = _RAND_48[20:0];
  _RAND_49 = {1{`RANDOM}};
  tag_regs_49 = _RAND_49[20:0];
  _RAND_50 = {1{`RANDOM}};
  tag_regs_50 = _RAND_50[20:0];
  _RAND_51 = {1{`RANDOM}};
  tag_regs_51 = _RAND_51[20:0];
  _RAND_52 = {1{`RANDOM}};
  tag_regs_52 = _RAND_52[20:0];
  _RAND_53 = {1{`RANDOM}};
  tag_regs_53 = _RAND_53[20:0];
  _RAND_54 = {1{`RANDOM}};
  tag_regs_54 = _RAND_54[20:0];
  _RAND_55 = {1{`RANDOM}};
  tag_regs_55 = _RAND_55[20:0];
  _RAND_56 = {1{`RANDOM}};
  tag_regs_56 = _RAND_56[20:0];
  _RAND_57 = {1{`RANDOM}};
  tag_regs_57 = _RAND_57[20:0];
  _RAND_58 = {1{`RANDOM}};
  tag_regs_58 = _RAND_58[20:0];
  _RAND_59 = {1{`RANDOM}};
  tag_regs_59 = _RAND_59[20:0];
  _RAND_60 = {1{`RANDOM}};
  tag_regs_60 = _RAND_60[20:0];
  _RAND_61 = {1{`RANDOM}};
  tag_regs_61 = _RAND_61[20:0];
  _RAND_62 = {1{`RANDOM}};
  tag_regs_62 = _RAND_62[20:0];
  _RAND_63 = {1{`RANDOM}};
  tag_regs_63 = _RAND_63[20:0];
  _RAND_64 = {1{`RANDOM}};
  tag_regs_64 = _RAND_64[20:0];
  _RAND_65 = {1{`RANDOM}};
  tag_regs_65 = _RAND_65[20:0];
  _RAND_66 = {1{`RANDOM}};
  tag_regs_66 = _RAND_66[20:0];
  _RAND_67 = {1{`RANDOM}};
  tag_regs_67 = _RAND_67[20:0];
  _RAND_68 = {1{`RANDOM}};
  tag_regs_68 = _RAND_68[20:0];
  _RAND_69 = {1{`RANDOM}};
  tag_regs_69 = _RAND_69[20:0];
  _RAND_70 = {1{`RANDOM}};
  tag_regs_70 = _RAND_70[20:0];
  _RAND_71 = {1{`RANDOM}};
  tag_regs_71 = _RAND_71[20:0];
  _RAND_72 = {1{`RANDOM}};
  tag_regs_72 = _RAND_72[20:0];
  _RAND_73 = {1{`RANDOM}};
  tag_regs_73 = _RAND_73[20:0];
  _RAND_74 = {1{`RANDOM}};
  tag_regs_74 = _RAND_74[20:0];
  _RAND_75 = {1{`RANDOM}};
  tag_regs_75 = _RAND_75[20:0];
  _RAND_76 = {1{`RANDOM}};
  tag_regs_76 = _RAND_76[20:0];
  _RAND_77 = {1{`RANDOM}};
  tag_regs_77 = _RAND_77[20:0];
  _RAND_78 = {1{`RANDOM}};
  tag_regs_78 = _RAND_78[20:0];
  _RAND_79 = {1{`RANDOM}};
  tag_regs_79 = _RAND_79[20:0];
  _RAND_80 = {1{`RANDOM}};
  tag_regs_80 = _RAND_80[20:0];
  _RAND_81 = {1{`RANDOM}};
  tag_regs_81 = _RAND_81[20:0];
  _RAND_82 = {1{`RANDOM}};
  tag_regs_82 = _RAND_82[20:0];
  _RAND_83 = {1{`RANDOM}};
  tag_regs_83 = _RAND_83[20:0];
  _RAND_84 = {1{`RANDOM}};
  tag_regs_84 = _RAND_84[20:0];
  _RAND_85 = {1{`RANDOM}};
  tag_regs_85 = _RAND_85[20:0];
  _RAND_86 = {1{`RANDOM}};
  tag_regs_86 = _RAND_86[20:0];
  _RAND_87 = {1{`RANDOM}};
  tag_regs_87 = _RAND_87[20:0];
  _RAND_88 = {1{`RANDOM}};
  tag_regs_88 = _RAND_88[20:0];
  _RAND_89 = {1{`RANDOM}};
  tag_regs_89 = _RAND_89[20:0];
  _RAND_90 = {1{`RANDOM}};
  tag_regs_90 = _RAND_90[20:0];
  _RAND_91 = {1{`RANDOM}};
  tag_regs_91 = _RAND_91[20:0];
  _RAND_92 = {1{`RANDOM}};
  tag_regs_92 = _RAND_92[20:0];
  _RAND_93 = {1{`RANDOM}};
  tag_regs_93 = _RAND_93[20:0];
  _RAND_94 = {1{`RANDOM}};
  tag_regs_94 = _RAND_94[20:0];
  _RAND_95 = {1{`RANDOM}};
  tag_regs_95 = _RAND_95[20:0];
  _RAND_96 = {1{`RANDOM}};
  tag_regs_96 = _RAND_96[20:0];
  _RAND_97 = {1{`RANDOM}};
  tag_regs_97 = _RAND_97[20:0];
  _RAND_98 = {1{`RANDOM}};
  tag_regs_98 = _RAND_98[20:0];
  _RAND_99 = {1{`RANDOM}};
  tag_regs_99 = _RAND_99[20:0];
  _RAND_100 = {1{`RANDOM}};
  tag_regs_100 = _RAND_100[20:0];
  _RAND_101 = {1{`RANDOM}};
  tag_regs_101 = _RAND_101[20:0];
  _RAND_102 = {1{`RANDOM}};
  tag_regs_102 = _RAND_102[20:0];
  _RAND_103 = {1{`RANDOM}};
  tag_regs_103 = _RAND_103[20:0];
  _RAND_104 = {1{`RANDOM}};
  tag_regs_104 = _RAND_104[20:0];
  _RAND_105 = {1{`RANDOM}};
  tag_regs_105 = _RAND_105[20:0];
  _RAND_106 = {1{`RANDOM}};
  tag_regs_106 = _RAND_106[20:0];
  _RAND_107 = {1{`RANDOM}};
  tag_regs_107 = _RAND_107[20:0];
  _RAND_108 = {1{`RANDOM}};
  tag_regs_108 = _RAND_108[20:0];
  _RAND_109 = {1{`RANDOM}};
  tag_regs_109 = _RAND_109[20:0];
  _RAND_110 = {1{`RANDOM}};
  tag_regs_110 = _RAND_110[20:0];
  _RAND_111 = {1{`RANDOM}};
  tag_regs_111 = _RAND_111[20:0];
  _RAND_112 = {1{`RANDOM}};
  tag_regs_112 = _RAND_112[20:0];
  _RAND_113 = {1{`RANDOM}};
  tag_regs_113 = _RAND_113[20:0];
  _RAND_114 = {1{`RANDOM}};
  tag_regs_114 = _RAND_114[20:0];
  _RAND_115 = {1{`RANDOM}};
  tag_regs_115 = _RAND_115[20:0];
  _RAND_116 = {1{`RANDOM}};
  tag_regs_116 = _RAND_116[20:0];
  _RAND_117 = {1{`RANDOM}};
  tag_regs_117 = _RAND_117[20:0];
  _RAND_118 = {1{`RANDOM}};
  tag_regs_118 = _RAND_118[20:0];
  _RAND_119 = {1{`RANDOM}};
  tag_regs_119 = _RAND_119[20:0];
  _RAND_120 = {1{`RANDOM}};
  tag_regs_120 = _RAND_120[20:0];
  _RAND_121 = {1{`RANDOM}};
  tag_regs_121 = _RAND_121[20:0];
  _RAND_122 = {1{`RANDOM}};
  tag_regs_122 = _RAND_122[20:0];
  _RAND_123 = {1{`RANDOM}};
  tag_regs_123 = _RAND_123[20:0];
  _RAND_124 = {1{`RANDOM}};
  tag_regs_124 = _RAND_124[20:0];
  _RAND_125 = {1{`RANDOM}};
  tag_regs_125 = _RAND_125[20:0];
  _RAND_126 = {1{`RANDOM}};
  tag_regs_126 = _RAND_126[20:0];
  _RAND_127 = {1{`RANDOM}};
  tag_regs_127 = _RAND_127[20:0];
  _RAND_128 = {1{`RANDOM}};
  tag_asid_regs_0 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  tag_asid_regs_1 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  tag_asid_regs_2 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  tag_asid_regs_3 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  tag_asid_regs_4 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  tag_asid_regs_5 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  tag_asid_regs_6 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  tag_asid_regs_7 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  tag_asid_regs_8 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  tag_asid_regs_9 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  tag_asid_regs_10 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  tag_asid_regs_11 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  tag_asid_regs_12 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  tag_asid_regs_13 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  tag_asid_regs_14 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  tag_asid_regs_15 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  tag_asid_regs_16 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  tag_asid_regs_17 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  tag_asid_regs_18 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  tag_asid_regs_19 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  tag_asid_regs_20 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  tag_asid_regs_21 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  tag_asid_regs_22 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  tag_asid_regs_23 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  tag_asid_regs_24 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  tag_asid_regs_25 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  tag_asid_regs_26 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  tag_asid_regs_27 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  tag_asid_regs_28 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  tag_asid_regs_29 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  tag_asid_regs_30 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  tag_asid_regs_31 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  tag_asid_regs_32 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  tag_asid_regs_33 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  tag_asid_regs_34 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  tag_asid_regs_35 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  tag_asid_regs_36 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  tag_asid_regs_37 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  tag_asid_regs_38 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  tag_asid_regs_39 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  tag_asid_regs_40 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  tag_asid_regs_41 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  tag_asid_regs_42 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  tag_asid_regs_43 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  tag_asid_regs_44 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  tag_asid_regs_45 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  tag_asid_regs_46 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  tag_asid_regs_47 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  tag_asid_regs_48 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  tag_asid_regs_49 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  tag_asid_regs_50 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  tag_asid_regs_51 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  tag_asid_regs_52 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  tag_asid_regs_53 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  tag_asid_regs_54 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  tag_asid_regs_55 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  tag_asid_regs_56 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  tag_asid_regs_57 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  tag_asid_regs_58 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  tag_asid_regs_59 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  tag_asid_regs_60 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  tag_asid_regs_61 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  tag_asid_regs_62 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  tag_asid_regs_63 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  tag_asid_regs_64 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  tag_asid_regs_65 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  tag_asid_regs_66 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  tag_asid_regs_67 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  tag_asid_regs_68 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  tag_asid_regs_69 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  tag_asid_regs_70 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  tag_asid_regs_71 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  tag_asid_regs_72 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  tag_asid_regs_73 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  tag_asid_regs_74 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  tag_asid_regs_75 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  tag_asid_regs_76 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  tag_asid_regs_77 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  tag_asid_regs_78 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  tag_asid_regs_79 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  tag_asid_regs_80 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  tag_asid_regs_81 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  tag_asid_regs_82 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  tag_asid_regs_83 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  tag_asid_regs_84 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  tag_asid_regs_85 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  tag_asid_regs_86 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  tag_asid_regs_87 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  tag_asid_regs_88 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  tag_asid_regs_89 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  tag_asid_regs_90 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  tag_asid_regs_91 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  tag_asid_regs_92 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  tag_asid_regs_93 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  tag_asid_regs_94 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  tag_asid_regs_95 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  tag_asid_regs_96 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  tag_asid_regs_97 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  tag_asid_regs_98 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  tag_asid_regs_99 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  tag_asid_regs_100 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  tag_asid_regs_101 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  tag_asid_regs_102 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  tag_asid_regs_103 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  tag_asid_regs_104 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  tag_asid_regs_105 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  tag_asid_regs_106 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  tag_asid_regs_107 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  tag_asid_regs_108 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  tag_asid_regs_109 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  tag_asid_regs_110 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  tag_asid_regs_111 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  tag_asid_regs_112 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  tag_asid_regs_113 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  tag_asid_regs_114 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  tag_asid_regs_115 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  tag_asid_regs_116 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  tag_asid_regs_117 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  tag_asid_regs_118 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  tag_asid_regs_119 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  tag_asid_regs_120 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  tag_asid_regs_121 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  tag_asid_regs_122 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  tag_asid_regs_123 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  tag_asid_regs_124 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  tag_asid_regs_125 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  tag_asid_regs_126 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  tag_asid_regs_127 = _RAND_255[7:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    tag_regs_0 = 21'h0;
  end
  if (reset) begin
    tag_regs_1 = 21'h0;
  end
  if (reset) begin
    tag_regs_2 = 21'h0;
  end
  if (reset) begin
    tag_regs_3 = 21'h0;
  end
  if (reset) begin
    tag_regs_4 = 21'h0;
  end
  if (reset) begin
    tag_regs_5 = 21'h0;
  end
  if (reset) begin
    tag_regs_6 = 21'h0;
  end
  if (reset) begin
    tag_regs_7 = 21'h0;
  end
  if (reset) begin
    tag_regs_8 = 21'h0;
  end
  if (reset) begin
    tag_regs_9 = 21'h0;
  end
  if (reset) begin
    tag_regs_10 = 21'h0;
  end
  if (reset) begin
    tag_regs_11 = 21'h0;
  end
  if (reset) begin
    tag_regs_12 = 21'h0;
  end
  if (reset) begin
    tag_regs_13 = 21'h0;
  end
  if (reset) begin
    tag_regs_14 = 21'h0;
  end
  if (reset) begin
    tag_regs_15 = 21'h0;
  end
  if (reset) begin
    tag_regs_16 = 21'h0;
  end
  if (reset) begin
    tag_regs_17 = 21'h0;
  end
  if (reset) begin
    tag_regs_18 = 21'h0;
  end
  if (reset) begin
    tag_regs_19 = 21'h0;
  end
  if (reset) begin
    tag_regs_20 = 21'h0;
  end
  if (reset) begin
    tag_regs_21 = 21'h0;
  end
  if (reset) begin
    tag_regs_22 = 21'h0;
  end
  if (reset) begin
    tag_regs_23 = 21'h0;
  end
  if (reset) begin
    tag_regs_24 = 21'h0;
  end
  if (reset) begin
    tag_regs_25 = 21'h0;
  end
  if (reset) begin
    tag_regs_26 = 21'h0;
  end
  if (reset) begin
    tag_regs_27 = 21'h0;
  end
  if (reset) begin
    tag_regs_28 = 21'h0;
  end
  if (reset) begin
    tag_regs_29 = 21'h0;
  end
  if (reset) begin
    tag_regs_30 = 21'h0;
  end
  if (reset) begin
    tag_regs_31 = 21'h0;
  end
  if (reset) begin
    tag_regs_32 = 21'h0;
  end
  if (reset) begin
    tag_regs_33 = 21'h0;
  end
  if (reset) begin
    tag_regs_34 = 21'h0;
  end
  if (reset) begin
    tag_regs_35 = 21'h0;
  end
  if (reset) begin
    tag_regs_36 = 21'h0;
  end
  if (reset) begin
    tag_regs_37 = 21'h0;
  end
  if (reset) begin
    tag_regs_38 = 21'h0;
  end
  if (reset) begin
    tag_regs_39 = 21'h0;
  end
  if (reset) begin
    tag_regs_40 = 21'h0;
  end
  if (reset) begin
    tag_regs_41 = 21'h0;
  end
  if (reset) begin
    tag_regs_42 = 21'h0;
  end
  if (reset) begin
    tag_regs_43 = 21'h0;
  end
  if (reset) begin
    tag_regs_44 = 21'h0;
  end
  if (reset) begin
    tag_regs_45 = 21'h0;
  end
  if (reset) begin
    tag_regs_46 = 21'h0;
  end
  if (reset) begin
    tag_regs_47 = 21'h0;
  end
  if (reset) begin
    tag_regs_48 = 21'h0;
  end
  if (reset) begin
    tag_regs_49 = 21'h0;
  end
  if (reset) begin
    tag_regs_50 = 21'h0;
  end
  if (reset) begin
    tag_regs_51 = 21'h0;
  end
  if (reset) begin
    tag_regs_52 = 21'h0;
  end
  if (reset) begin
    tag_regs_53 = 21'h0;
  end
  if (reset) begin
    tag_regs_54 = 21'h0;
  end
  if (reset) begin
    tag_regs_55 = 21'h0;
  end
  if (reset) begin
    tag_regs_56 = 21'h0;
  end
  if (reset) begin
    tag_regs_57 = 21'h0;
  end
  if (reset) begin
    tag_regs_58 = 21'h0;
  end
  if (reset) begin
    tag_regs_59 = 21'h0;
  end
  if (reset) begin
    tag_regs_60 = 21'h0;
  end
  if (reset) begin
    tag_regs_61 = 21'h0;
  end
  if (reset) begin
    tag_regs_62 = 21'h0;
  end
  if (reset) begin
    tag_regs_63 = 21'h0;
  end
  if (reset) begin
    tag_regs_64 = 21'h0;
  end
  if (reset) begin
    tag_regs_65 = 21'h0;
  end
  if (reset) begin
    tag_regs_66 = 21'h0;
  end
  if (reset) begin
    tag_regs_67 = 21'h0;
  end
  if (reset) begin
    tag_regs_68 = 21'h0;
  end
  if (reset) begin
    tag_regs_69 = 21'h0;
  end
  if (reset) begin
    tag_regs_70 = 21'h0;
  end
  if (reset) begin
    tag_regs_71 = 21'h0;
  end
  if (reset) begin
    tag_regs_72 = 21'h0;
  end
  if (reset) begin
    tag_regs_73 = 21'h0;
  end
  if (reset) begin
    tag_regs_74 = 21'h0;
  end
  if (reset) begin
    tag_regs_75 = 21'h0;
  end
  if (reset) begin
    tag_regs_76 = 21'h0;
  end
  if (reset) begin
    tag_regs_77 = 21'h0;
  end
  if (reset) begin
    tag_regs_78 = 21'h0;
  end
  if (reset) begin
    tag_regs_79 = 21'h0;
  end
  if (reset) begin
    tag_regs_80 = 21'h0;
  end
  if (reset) begin
    tag_regs_81 = 21'h0;
  end
  if (reset) begin
    tag_regs_82 = 21'h0;
  end
  if (reset) begin
    tag_regs_83 = 21'h0;
  end
  if (reset) begin
    tag_regs_84 = 21'h0;
  end
  if (reset) begin
    tag_regs_85 = 21'h0;
  end
  if (reset) begin
    tag_regs_86 = 21'h0;
  end
  if (reset) begin
    tag_regs_87 = 21'h0;
  end
  if (reset) begin
    tag_regs_88 = 21'h0;
  end
  if (reset) begin
    tag_regs_89 = 21'h0;
  end
  if (reset) begin
    tag_regs_90 = 21'h0;
  end
  if (reset) begin
    tag_regs_91 = 21'h0;
  end
  if (reset) begin
    tag_regs_92 = 21'h0;
  end
  if (reset) begin
    tag_regs_93 = 21'h0;
  end
  if (reset) begin
    tag_regs_94 = 21'h0;
  end
  if (reset) begin
    tag_regs_95 = 21'h0;
  end
  if (reset) begin
    tag_regs_96 = 21'h0;
  end
  if (reset) begin
    tag_regs_97 = 21'h0;
  end
  if (reset) begin
    tag_regs_98 = 21'h0;
  end
  if (reset) begin
    tag_regs_99 = 21'h0;
  end
  if (reset) begin
    tag_regs_100 = 21'h0;
  end
  if (reset) begin
    tag_regs_101 = 21'h0;
  end
  if (reset) begin
    tag_regs_102 = 21'h0;
  end
  if (reset) begin
    tag_regs_103 = 21'h0;
  end
  if (reset) begin
    tag_regs_104 = 21'h0;
  end
  if (reset) begin
    tag_regs_105 = 21'h0;
  end
  if (reset) begin
    tag_regs_106 = 21'h0;
  end
  if (reset) begin
    tag_regs_107 = 21'h0;
  end
  if (reset) begin
    tag_regs_108 = 21'h0;
  end
  if (reset) begin
    tag_regs_109 = 21'h0;
  end
  if (reset) begin
    tag_regs_110 = 21'h0;
  end
  if (reset) begin
    tag_regs_111 = 21'h0;
  end
  if (reset) begin
    tag_regs_112 = 21'h0;
  end
  if (reset) begin
    tag_regs_113 = 21'h0;
  end
  if (reset) begin
    tag_regs_114 = 21'h0;
  end
  if (reset) begin
    tag_regs_115 = 21'h0;
  end
  if (reset) begin
    tag_regs_116 = 21'h0;
  end
  if (reset) begin
    tag_regs_117 = 21'h0;
  end
  if (reset) begin
    tag_regs_118 = 21'h0;
  end
  if (reset) begin
    tag_regs_119 = 21'h0;
  end
  if (reset) begin
    tag_regs_120 = 21'h0;
  end
  if (reset) begin
    tag_regs_121 = 21'h0;
  end
  if (reset) begin
    tag_regs_122 = 21'h0;
  end
  if (reset) begin
    tag_regs_123 = 21'h0;
  end
  if (reset) begin
    tag_regs_124 = 21'h0;
  end
  if (reset) begin
    tag_regs_125 = 21'h0;
  end
  if (reset) begin
    tag_regs_126 = 21'h0;
  end
  if (reset) begin
    tag_regs_127 = 21'h0;
  end
  if (reset) begin
    tag_asid_regs_0 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_1 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_2 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_3 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_4 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_5 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_6 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_7 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_8 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_9 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_10 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_11 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_12 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_13 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_14 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_15 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_16 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_17 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_18 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_19 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_20 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_21 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_22 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_23 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_24 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_25 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_26 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_27 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_28 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_29 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_30 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_31 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_32 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_33 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_34 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_35 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_36 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_37 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_38 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_39 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_40 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_41 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_42 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_43 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_44 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_45 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_46 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_47 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_48 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_49 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_50 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_51 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_52 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_53 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_54 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_55 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_56 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_57 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_58 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_59 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_60 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_61 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_62 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_63 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_64 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_65 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_66 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_67 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_68 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_69 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_70 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_71 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_72 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_73 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_74 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_75 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_76 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_77 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_78 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_79 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_80 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_81 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_82 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_83 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_84 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_85 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_86 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_87 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_88 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_89 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_90 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_91 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_92 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_93 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_94 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_95 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_96 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_97 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_98 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_99 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_100 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_101 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_102 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_103 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_104 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_105 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_106 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_107 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_108 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_109 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_110 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_111 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_112 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_113 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_114 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_115 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_116 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_117 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_118 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_119 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_120 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_121 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_122 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_123 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_124 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_125 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_126 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_127 = 8'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module icache_data(
  input         clock,
  input  [4:0]  io_wen,
  input  [31:0] io_addr,
  input  [39:0] io_wdata,
  output [39:0] io_rdata
);
  wire  icache_data_ram_0_clka; // @[icache_data.scala 32:35]
  wire  icache_data_ram_0_ena; // @[icache_data.scala 32:35]
  wire [4:0] icache_data_ram_0_wea; // @[icache_data.scala 32:35]
  wire [6:0] icache_data_ram_0_addra; // @[icache_data.scala 32:35]
  wire [39:0] icache_data_ram_0_dina; // @[icache_data.scala 32:35]
  wire [39:0] icache_data_ram_0_douta; // @[icache_data.scala 32:35]
  icache_data_ram icache_data_ram_0 ( // @[icache_data.scala 32:35]
    .clka(icache_data_ram_0_clka),
    .ena(icache_data_ram_0_ena),
    .wea(icache_data_ram_0_wea),
    .addra(icache_data_ram_0_addra),
    .dina(icache_data_ram_0_dina),
    .douta(icache_data_ram_0_douta)
  );
  assign io_rdata = icache_data_ram_0_douta; // @[icache_data.scala 38:18]
  assign icache_data_ram_0_clka = clock; // @[icache_data.scala 33:40]
  assign icache_data_ram_0_ena = 1'h1; // @[icache_data.scala 34:32]
  assign icache_data_ram_0_wea = io_wen; // @[icache_data.scala 35:31]
  assign icache_data_ram_0_addra = io_addr[11:5]; // @[icache_data.scala 36:42]
  assign icache_data_ram_0_dina = io_wdata; // @[icache_data.scala 37:31]
endmodule
module inst_cache(
  input         clock,
  input         reset,
  output [31:0] io_port_araddr,
  output [3:0]  io_port_arlen,
  output [1:0]  io_port_arburst,
  output        io_port_arvalid,
  input         io_port_arready,
  input  [31:0] io_port_rdata,
  input         io_port_rlast,
  input         io_port_rvalid,
  input         io_port_sram_req,
  input  [31:0] io_port_sram_addr,
  output [1:0]  io_port_sram_write_en,
  output [39:0] io_port_sram_rdata_L,
  input         io_port_sram_cache,
  input         io_stage2_flush,
  output        io_stage2_stall,
  input  [1:0]  io_stage1_valid_flush,
  input         io_inst_ready_to_use,
  input         io_inst_buffer_full,
  output [1:0]  io_stage2_exception,
  input  [7:0]  io_cp0_asid,
  output [31:0] io_v_addr_for_tlb,
  input  [31:0] io_p_addr_for_tlb,
  output        io_tlb_req,
  input  [1:0]  io_tlb_exception,
  input         io_inst_ready_branch,
  input         io_inst_buffer_empty
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [63:0] _RAND_145;
`endif // RANDOMIZE_REG_INIT
  wire  icache_tag_clock; // @[inst_cache.scala 93:34]
  wire  icache_tag_reset; // @[inst_cache.scala 93:34]
  wire  icache_tag_io_wen; // @[inst_cache.scala 93:34]
  wire [20:0] icache_tag_io_wdata; // @[inst_cache.scala 93:34]
  wire [31:0] icache_tag_io_addr; // @[inst_cache.scala 93:34]
  wire  icache_tag_io_hit; // @[inst_cache.scala 93:34]
  wire  icache_tag_io_valid; // @[inst_cache.scala 93:34]
  wire [7:0] icache_tag_io_asid; // @[inst_cache.scala 93:34]
  wire  icache_tag_1_clock; // @[inst_cache.scala 95:34]
  wire  icache_tag_1_reset; // @[inst_cache.scala 95:34]
  wire  icache_tag_1_io_wen; // @[inst_cache.scala 95:34]
  wire [20:0] icache_tag_1_io_wdata; // @[inst_cache.scala 95:34]
  wire [31:0] icache_tag_1_io_addr; // @[inst_cache.scala 95:34]
  wire  icache_tag_1_io_hit; // @[inst_cache.scala 95:34]
  wire  icache_tag_1_io_valid; // @[inst_cache.scala 95:34]
  wire [7:0] icache_tag_1_io_asid; // @[inst_cache.scala 95:34]
  wire  icache_data_clock; // @[inst_cache.scala 98:55]
  wire [4:0] icache_data_io_wen; // @[inst_cache.scala 98:55]
  wire [31:0] icache_data_io_addr; // @[inst_cache.scala 98:55]
  wire [39:0] icache_data_io_wdata; // @[inst_cache.scala 98:55]
  wire [39:0] icache_data_io_rdata; // @[inst_cache.scala 98:55]
  wire  icache_data_1_clock; // @[inst_cache.scala 98:55]
  wire [4:0] icache_data_1_io_wen; // @[inst_cache.scala 98:55]
  wire [31:0] icache_data_1_io_addr; // @[inst_cache.scala 98:55]
  wire [39:0] icache_data_1_io_wdata; // @[inst_cache.scala 98:55]
  wire [39:0] icache_data_1_io_rdata; // @[inst_cache.scala 98:55]
  wire  icache_data_2_clock; // @[inst_cache.scala 98:55]
  wire [4:0] icache_data_2_io_wen; // @[inst_cache.scala 98:55]
  wire [31:0] icache_data_2_io_addr; // @[inst_cache.scala 98:55]
  wire [39:0] icache_data_2_io_wdata; // @[inst_cache.scala 98:55]
  wire [39:0] icache_data_2_io_rdata; // @[inst_cache.scala 98:55]
  wire  icache_data_3_clock; // @[inst_cache.scala 98:55]
  wire [4:0] icache_data_3_io_wen; // @[inst_cache.scala 98:55]
  wire [31:0] icache_data_3_io_addr; // @[inst_cache.scala 98:55]
  wire [39:0] icache_data_3_io_wdata; // @[inst_cache.scala 98:55]
  wire [39:0] icache_data_3_io_rdata; // @[inst_cache.scala 98:55]
  wire  icache_data_4_clock; // @[inst_cache.scala 98:55]
  wire [4:0] icache_data_4_io_wen; // @[inst_cache.scala 98:55]
  wire [31:0] icache_data_4_io_addr; // @[inst_cache.scala 98:55]
  wire [39:0] icache_data_4_io_wdata; // @[inst_cache.scala 98:55]
  wire [39:0] icache_data_4_io_rdata; // @[inst_cache.scala 98:55]
  wire  icache_data_5_clock; // @[inst_cache.scala 98:55]
  wire [4:0] icache_data_5_io_wen; // @[inst_cache.scala 98:55]
  wire [31:0] icache_data_5_io_addr; // @[inst_cache.scala 98:55]
  wire [39:0] icache_data_5_io_wdata; // @[inst_cache.scala 98:55]
  wire [39:0] icache_data_5_io_rdata; // @[inst_cache.scala 98:55]
  wire  icache_data_6_clock; // @[inst_cache.scala 98:55]
  wire [4:0] icache_data_6_io_wen; // @[inst_cache.scala 98:55]
  wire [31:0] icache_data_6_io_addr; // @[inst_cache.scala 98:55]
  wire [39:0] icache_data_6_io_wdata; // @[inst_cache.scala 98:55]
  wire [39:0] icache_data_6_io_rdata; // @[inst_cache.scala 98:55]
  wire  icache_data_7_clock; // @[inst_cache.scala 98:55]
  wire [4:0] icache_data_7_io_wen; // @[inst_cache.scala 98:55]
  wire [31:0] icache_data_7_io_addr; // @[inst_cache.scala 98:55]
  wire [39:0] icache_data_7_io_wdata; // @[inst_cache.scala 98:55]
  wire [39:0] icache_data_7_io_rdata; // @[inst_cache.scala 98:55]
  wire  icache_data_8_clock; // @[inst_cache.scala 99:55]
  wire [4:0] icache_data_8_io_wen; // @[inst_cache.scala 99:55]
  wire [31:0] icache_data_8_io_addr; // @[inst_cache.scala 99:55]
  wire [39:0] icache_data_8_io_wdata; // @[inst_cache.scala 99:55]
  wire [39:0] icache_data_8_io_rdata; // @[inst_cache.scala 99:55]
  wire  icache_data_9_clock; // @[inst_cache.scala 99:55]
  wire [4:0] icache_data_9_io_wen; // @[inst_cache.scala 99:55]
  wire [31:0] icache_data_9_io_addr; // @[inst_cache.scala 99:55]
  wire [39:0] icache_data_9_io_wdata; // @[inst_cache.scala 99:55]
  wire [39:0] icache_data_9_io_rdata; // @[inst_cache.scala 99:55]
  wire  icache_data_10_clock; // @[inst_cache.scala 99:55]
  wire [4:0] icache_data_10_io_wen; // @[inst_cache.scala 99:55]
  wire [31:0] icache_data_10_io_addr; // @[inst_cache.scala 99:55]
  wire [39:0] icache_data_10_io_wdata; // @[inst_cache.scala 99:55]
  wire [39:0] icache_data_10_io_rdata; // @[inst_cache.scala 99:55]
  wire  icache_data_11_clock; // @[inst_cache.scala 99:55]
  wire [4:0] icache_data_11_io_wen; // @[inst_cache.scala 99:55]
  wire [31:0] icache_data_11_io_addr; // @[inst_cache.scala 99:55]
  wire [39:0] icache_data_11_io_wdata; // @[inst_cache.scala 99:55]
  wire [39:0] icache_data_11_io_rdata; // @[inst_cache.scala 99:55]
  wire  icache_data_12_clock; // @[inst_cache.scala 99:55]
  wire [4:0] icache_data_12_io_wen; // @[inst_cache.scala 99:55]
  wire [31:0] icache_data_12_io_addr; // @[inst_cache.scala 99:55]
  wire [39:0] icache_data_12_io_wdata; // @[inst_cache.scala 99:55]
  wire [39:0] icache_data_12_io_rdata; // @[inst_cache.scala 99:55]
  wire  icache_data_13_clock; // @[inst_cache.scala 99:55]
  wire [4:0] icache_data_13_io_wen; // @[inst_cache.scala 99:55]
  wire [31:0] icache_data_13_io_addr; // @[inst_cache.scala 99:55]
  wire [39:0] icache_data_13_io_wdata; // @[inst_cache.scala 99:55]
  wire [39:0] icache_data_13_io_rdata; // @[inst_cache.scala 99:55]
  wire  icache_data_14_clock; // @[inst_cache.scala 99:55]
  wire [4:0] icache_data_14_io_wen; // @[inst_cache.scala 99:55]
  wire [31:0] icache_data_14_io_addr; // @[inst_cache.scala 99:55]
  wire [39:0] icache_data_14_io_wdata; // @[inst_cache.scala 99:55]
  wire [39:0] icache_data_14_io_rdata; // @[inst_cache.scala 99:55]
  wire  icache_data_15_clock; // @[inst_cache.scala 99:55]
  wire [4:0] icache_data_15_io_wen; // @[inst_cache.scala 99:55]
  wire [31:0] icache_data_15_io_addr; // @[inst_cache.scala 99:55]
  wire [39:0] icache_data_15_io_wdata; // @[inst_cache.scala 99:55]
  wire [39:0] icache_data_15_io_rdata; // @[inst_cache.scala 99:55]
  reg  lru_0; // @[inst_cache.scala 86:22]
  reg  lru_1; // @[inst_cache.scala 86:22]
  reg  lru_2; // @[inst_cache.scala 86:22]
  reg  lru_3; // @[inst_cache.scala 86:22]
  reg  lru_4; // @[inst_cache.scala 86:22]
  reg  lru_5; // @[inst_cache.scala 86:22]
  reg  lru_6; // @[inst_cache.scala 86:22]
  reg  lru_7; // @[inst_cache.scala 86:22]
  reg  lru_8; // @[inst_cache.scala 86:22]
  reg  lru_9; // @[inst_cache.scala 86:22]
  reg  lru_10; // @[inst_cache.scala 86:22]
  reg  lru_11; // @[inst_cache.scala 86:22]
  reg  lru_12; // @[inst_cache.scala 86:22]
  reg  lru_13; // @[inst_cache.scala 86:22]
  reg  lru_14; // @[inst_cache.scala 86:22]
  reg  lru_15; // @[inst_cache.scala 86:22]
  reg  lru_16; // @[inst_cache.scala 86:22]
  reg  lru_17; // @[inst_cache.scala 86:22]
  reg  lru_18; // @[inst_cache.scala 86:22]
  reg  lru_19; // @[inst_cache.scala 86:22]
  reg  lru_20; // @[inst_cache.scala 86:22]
  reg  lru_21; // @[inst_cache.scala 86:22]
  reg  lru_22; // @[inst_cache.scala 86:22]
  reg  lru_23; // @[inst_cache.scala 86:22]
  reg  lru_24; // @[inst_cache.scala 86:22]
  reg  lru_25; // @[inst_cache.scala 86:22]
  reg  lru_26; // @[inst_cache.scala 86:22]
  reg  lru_27; // @[inst_cache.scala 86:22]
  reg  lru_28; // @[inst_cache.scala 86:22]
  reg  lru_29; // @[inst_cache.scala 86:22]
  reg  lru_30; // @[inst_cache.scala 86:22]
  reg  lru_31; // @[inst_cache.scala 86:22]
  reg  lru_32; // @[inst_cache.scala 86:22]
  reg  lru_33; // @[inst_cache.scala 86:22]
  reg  lru_34; // @[inst_cache.scala 86:22]
  reg  lru_35; // @[inst_cache.scala 86:22]
  reg  lru_36; // @[inst_cache.scala 86:22]
  reg  lru_37; // @[inst_cache.scala 86:22]
  reg  lru_38; // @[inst_cache.scala 86:22]
  reg  lru_39; // @[inst_cache.scala 86:22]
  reg  lru_40; // @[inst_cache.scala 86:22]
  reg  lru_41; // @[inst_cache.scala 86:22]
  reg  lru_42; // @[inst_cache.scala 86:22]
  reg  lru_43; // @[inst_cache.scala 86:22]
  reg  lru_44; // @[inst_cache.scala 86:22]
  reg  lru_45; // @[inst_cache.scala 86:22]
  reg  lru_46; // @[inst_cache.scala 86:22]
  reg  lru_47; // @[inst_cache.scala 86:22]
  reg  lru_48; // @[inst_cache.scala 86:22]
  reg  lru_49; // @[inst_cache.scala 86:22]
  reg  lru_50; // @[inst_cache.scala 86:22]
  reg  lru_51; // @[inst_cache.scala 86:22]
  reg  lru_52; // @[inst_cache.scala 86:22]
  reg  lru_53; // @[inst_cache.scala 86:22]
  reg  lru_54; // @[inst_cache.scala 86:22]
  reg  lru_55; // @[inst_cache.scala 86:22]
  reg  lru_56; // @[inst_cache.scala 86:22]
  reg  lru_57; // @[inst_cache.scala 86:22]
  reg  lru_58; // @[inst_cache.scala 86:22]
  reg  lru_59; // @[inst_cache.scala 86:22]
  reg  lru_60; // @[inst_cache.scala 86:22]
  reg  lru_61; // @[inst_cache.scala 86:22]
  reg  lru_62; // @[inst_cache.scala 86:22]
  reg  lru_63; // @[inst_cache.scala 86:22]
  reg  lru_64; // @[inst_cache.scala 86:22]
  reg  lru_65; // @[inst_cache.scala 86:22]
  reg  lru_66; // @[inst_cache.scala 86:22]
  reg  lru_67; // @[inst_cache.scala 86:22]
  reg  lru_68; // @[inst_cache.scala 86:22]
  reg  lru_69; // @[inst_cache.scala 86:22]
  reg  lru_70; // @[inst_cache.scala 86:22]
  reg  lru_71; // @[inst_cache.scala 86:22]
  reg  lru_72; // @[inst_cache.scala 86:22]
  reg  lru_73; // @[inst_cache.scala 86:22]
  reg  lru_74; // @[inst_cache.scala 86:22]
  reg  lru_75; // @[inst_cache.scala 86:22]
  reg  lru_76; // @[inst_cache.scala 86:22]
  reg  lru_77; // @[inst_cache.scala 86:22]
  reg  lru_78; // @[inst_cache.scala 86:22]
  reg  lru_79; // @[inst_cache.scala 86:22]
  reg  lru_80; // @[inst_cache.scala 86:22]
  reg  lru_81; // @[inst_cache.scala 86:22]
  reg  lru_82; // @[inst_cache.scala 86:22]
  reg  lru_83; // @[inst_cache.scala 86:22]
  reg  lru_84; // @[inst_cache.scala 86:22]
  reg  lru_85; // @[inst_cache.scala 86:22]
  reg  lru_86; // @[inst_cache.scala 86:22]
  reg  lru_87; // @[inst_cache.scala 86:22]
  reg  lru_88; // @[inst_cache.scala 86:22]
  reg  lru_89; // @[inst_cache.scala 86:22]
  reg  lru_90; // @[inst_cache.scala 86:22]
  reg  lru_91; // @[inst_cache.scala 86:22]
  reg  lru_92; // @[inst_cache.scala 86:22]
  reg  lru_93; // @[inst_cache.scala 86:22]
  reg  lru_94; // @[inst_cache.scala 86:22]
  reg  lru_95; // @[inst_cache.scala 86:22]
  reg  lru_96; // @[inst_cache.scala 86:22]
  reg  lru_97; // @[inst_cache.scala 86:22]
  reg  lru_98; // @[inst_cache.scala 86:22]
  reg  lru_99; // @[inst_cache.scala 86:22]
  reg  lru_100; // @[inst_cache.scala 86:22]
  reg  lru_101; // @[inst_cache.scala 86:22]
  reg  lru_102; // @[inst_cache.scala 86:22]
  reg  lru_103; // @[inst_cache.scala 86:22]
  reg  lru_104; // @[inst_cache.scala 86:22]
  reg  lru_105; // @[inst_cache.scala 86:22]
  reg  lru_106; // @[inst_cache.scala 86:22]
  reg  lru_107; // @[inst_cache.scala 86:22]
  reg  lru_108; // @[inst_cache.scala 86:22]
  reg  lru_109; // @[inst_cache.scala 86:22]
  reg  lru_110; // @[inst_cache.scala 86:22]
  reg  lru_111; // @[inst_cache.scala 86:22]
  reg  lru_112; // @[inst_cache.scala 86:22]
  reg  lru_113; // @[inst_cache.scala 86:22]
  reg  lru_114; // @[inst_cache.scala 86:22]
  reg  lru_115; // @[inst_cache.scala 86:22]
  reg  lru_116; // @[inst_cache.scala 86:22]
  reg  lru_117; // @[inst_cache.scala 86:22]
  reg  lru_118; // @[inst_cache.scala 86:22]
  reg  lru_119; // @[inst_cache.scala 86:22]
  reg  lru_120; // @[inst_cache.scala 86:22]
  reg  lru_121; // @[inst_cache.scala 86:22]
  reg  lru_122; // @[inst_cache.scala 86:22]
  reg  lru_123; // @[inst_cache.scala 86:22]
  reg  lru_124; // @[inst_cache.scala 86:22]
  reg  lru_125; // @[inst_cache.scala 86:22]
  reg  lru_126; // @[inst_cache.scala 86:22]
  reg  lru_127; // @[inst_cache.scala 86:22]
  reg [3:0] work_state; // @[inst_cache.scala 110:29]
  reg [2:0] write_counter; // @[inst_cache.scala 112:33]
  reg [39:0] wait_data_L; // @[inst_cache.scala 113:31]
  reg  stage1_stall_reg; // @[inst_cache.scala 126:35]
  reg [31:0] stage1_sram_addr_reg; // @[Reg.scala 28:20]
  reg [31:0] stage1_sram_phy_addr_reg; // @[inst_cache.scala 130:43]
  reg  stage1_sram_cache_reg; // @[Reg.scala 28:20]
  reg  stage1_sram_req_reg; // @[Reg.scala 28:20]
  reg [1:0] stage1_sram_valid; // @[inst_cache.scala 133:36]
  reg  stage1_finished; // @[inst_cache.scala 135:34]
  reg [1:0] stage1_exception; // @[inst_cache.scala 136:35]
  reg [1:0] stage2_exception; // @[inst_cache.scala 140:35]
  wire [31:0] _stage1_sram_phy_addr_reg_T = io_tlb_req ? io_p_addr_for_tlb : stage1_sram_addr_reg; // @[inst_cache.scala 146:74]
  wire [31:0] _stage1_sram_phy_addr_reg_T_4 = {3'h0,_stage1_sram_phy_addr_reg_T[28:0]}; // @[Cat.scala 31:58]
  wire  _stage1_finished_T_1 = work_state == 4'h7; // @[inst_cache.scala 152:67]
  wire  _stage1_finished_T_2 = work_state == 4'h3; // @[inst_cache.scala 152:103]
  wire [1:0] _access_stage1_sram_valid_T_2 = io_stage1_valid_flush[1] ? 2'h2 : stage1_sram_valid; // @[inst_cache.scala 154:12]
  wire [1:0] access_stage1_sram_valid = io_stage1_valid_flush[0] ? 2'h1 : _access_stage1_sram_valid_T_2; // @[inst_cache.scala 153:40]
  wire  _access_work_state_T = work_state == 4'h2; // @[inst_cache.scala 256:41]
  wire  _access_work_state_T_6 = io_port_rlast & io_port_rvalid; // @[inst_cache.scala 257:71]
  wire [2:0] _access_work_state_T_7 = io_port_rlast & io_port_rvalid ? 3'h4 : 3'h3; // @[inst_cache.scala 257:49]
  wire  _access_work_state_T_8 = work_state == 4'h4; // @[inst_cache.scala 258:23]
  wire  _hit_T = icache_tag_io_hit; // @[inst_cache.scala 182:33]
  wire  _hit_T_2 = icache_tag_io_hit & icache_tag_io_valid; // @[inst_cache.scala 182:40]
  wire  _hit_T_3 = icache_tag_1_io_hit; // @[inst_cache.scala 183:27]
  wire  _hit_T_5 = icache_tag_1_io_hit & icache_tag_1_io_valid; // @[inst_cache.scala 183:34]
  wire  hit = icache_tag_io_hit & icache_tag_io_valid | _hit_T_5; // @[inst_cache.scala 182:70]
  wire [2:0] _access_work_state_T_13 = stage1_finished ? 3'h4 : 3'h2; // @[inst_cache.scala 258:145]
  wire [2:0] _access_work_state_T_14 = stage1_sram_cache_reg ? 3'h1 : _access_work_state_T_13; // @[inst_cache.scala 258:99]
  wire [2:0] _access_work_state_T_15 = stage1_sram_req_reg ? _access_work_state_T_14 : 3'h1; // @[inst_cache.scala 258:68]
  wire [2:0] _access_work_state_T_18 = stage1_finished ? 3'h4 : 3'h5; // @[inst_cache.scala 259:79]
  wire [2:0] _access_work_state_T_20 = stage1_sram_cache_reg ? _access_work_state_T_18 : _access_work_state_T_13; // @[inst_cache.scala 259:46]
  wire [2:0] _access_work_state_T_21 = stage1_sram_req_reg ? _access_work_state_T_20 : 3'h1; // @[inst_cache.scala 259:15]
  wire [2:0] _access_work_state_T_22 = hit ? _access_work_state_T_15 : _access_work_state_T_21; // @[inst_cache.scala 258:46]
  wire  _access_work_state_T_23 = work_state == 4'h1; // @[inst_cache.scala 261:23]
  wire [1:0] _access_work_state_T_28 = stage1_sram_cache_reg ? 2'h1 : 2'h2; // @[inst_cache.scala 261:95]
  wire [1:0] _access_work_state_T_29 = stage1_sram_req_reg ? _access_work_state_T_28 : 2'h1; // @[inst_cache.scala 261:64]
  wire [2:0] _access_work_state_T_32 = stage1_sram_cache_reg ? 3'h5 : 3'h2; // @[inst_cache.scala 262:46]
  wire [2:0] _access_work_state_T_33 = stage1_sram_req_reg ? _access_work_state_T_32 : 3'h1; // @[inst_cache.scala 262:15]
  wire [2:0] _access_work_state_T_34 = hit ? {{1'd0}, _access_work_state_T_29} : _access_work_state_T_33; // @[inst_cache.scala 261:42]
  wire  _access_work_state_T_35 = work_state == 4'h5; // @[inst_cache.scala 263:23]
  wire  _access_work_state_T_38 = work_state == 4'h6; // @[inst_cache.scala 264:23]
  wire [3:0] _access_work_state_T_42 = _access_work_state_T_6 ? 4'h7 : work_state; // @[inst_cache.scala 264:54]
  wire [3:0] _access_work_state_T_44 = _stage1_finished_T_1 ? 4'h4 : work_state; // @[inst_cache.scala 265:12]
  wire [3:0] _access_work_state_T_45 = work_state == 4'h6 ? _access_work_state_T_42 : _access_work_state_T_44; // @[inst_cache.scala 264:12]
  wire [3:0] _access_work_state_T_46 = work_state == 4'h5 & io_port_arready ? 4'h6 : _access_work_state_T_45; // @[inst_cache.scala 263:12]
  wire [3:0] _access_work_state_T_47 = work_state == 4'h1 ? {{1'd0}, _access_work_state_T_34} : _access_work_state_T_46; // @[inst_cache.scala 261:12]
  wire [3:0] _access_work_state_T_48 = work_state == 4'h4 ? {{1'd0}, _access_work_state_T_22} : _access_work_state_T_47; // @[inst_cache.scala 258:12]
  wire [3:0] _access_work_state_T_49 = _stage1_finished_T_2 ? {{1'd0}, _access_work_state_T_7} : _access_work_state_T_48
    ; // @[inst_cache.scala 257:12]
  wire [3:0] access_work_state = work_state == 4'h2 & io_port_arready ? 4'h3 : _access_work_state_T_49; // @[inst_cache.scala 256:30]
  wire  _stage2_stall_T = access_work_state == 4'h1; // @[inst_cache.scala 156:40]
  wire  _stage2_stall_T_3 = stage1_exception != 2'h0; // @[inst_cache.scala 156:120]
  wire  _stage2_stall_T_5 = ~io_inst_buffer_full; // @[inst_cache.scala 157:11]
  wire  stage2_stall = (access_work_state == 4'h1 | access_work_state == 4'h4 | stage1_exception != 2'h0) &
    _stage2_stall_T_5; // @[inst_cache.scala 156:129]
  wire [5:0] decoder_inst_data_opD = io_port_rdata[31:26]; // @[inst_cache.scala 69:24]
  wire [4:0] decoder_inst_data_RtD = io_port_rdata[20:16]; // @[inst_cache.scala 70:24]
  wire [5:0] decoder_inst_data_FunctD = io_port_rdata[5:0]; // @[inst_cache.scala 71:27]
  wire [2:0] _decoder_inst_data_T_1 = 5'h1 == decoder_inst_data_RtD ? 3'h4 : 3'h0; // @[Mux.scala 81:58]
  wire [2:0] _decoder_inst_data_T_3 = 5'h11 == decoder_inst_data_RtD ? 3'h4 : _decoder_inst_data_T_1; // @[Mux.scala 81:58]
  wire [5:0] _decoder_inst_data_T_5 = 5'h0 == decoder_inst_data_RtD ? 6'h20 : {{3'd0}, _decoder_inst_data_T_3}; // @[Mux.scala 81:58]
  wire [5:0] _decoder_inst_data_T_7 = 5'h10 == decoder_inst_data_RtD ? 6'h20 : _decoder_inst_data_T_5; // @[Mux.scala 81:58]
  wire [1:0] _decoder_inst_data_T_11 = 6'h5 == decoder_inst_data_opD ? 2'h2 : {{1'd0}, 6'h4 == decoder_inst_data_opD}; // @[Mux.scala 81:58]
  wire [3:0] _decoder_inst_data_T_13 = 6'h7 == decoder_inst_data_opD ? 4'h8 : {{2'd0}, _decoder_inst_data_T_11}; // @[Mux.scala 81:58]
  wire [4:0] _decoder_inst_data_T_15 = 6'h6 == decoder_inst_data_opD ? 5'h10 : {{1'd0}, _decoder_inst_data_T_13}; // @[Mux.scala 81:58]
  wire [5:0] _decoder_inst_data_T_17 = 6'h1 == decoder_inst_data_opD ? _decoder_inst_data_T_7 : {{1'd0},
    _decoder_inst_data_T_15}; // @[Mux.scala 81:58]
  wire  _decoder_inst_data_T_27 = 6'h0 == decoder_inst_data_opD ? 6'h9 == decoder_inst_data_FunctD | 6'h8 ==
    decoder_inst_data_FunctD : 6'h3 == decoder_inst_data_opD | 6'h2 == decoder_inst_data_opD; // @[Mux.scala 81:58]
  wire  _decoder_inst_data_T_45 = 6'h1 == decoder_inst_data_opD ? 5'h10 == decoder_inst_data_RtD | (5'h0 ==
    decoder_inst_data_RtD | (5'h11 == decoder_inst_data_RtD | 5'h1 == decoder_inst_data_RtD)) : 6'h6 ==
    decoder_inst_data_opD | (6'h7 == decoder_inst_data_opD | (6'h5 == decoder_inst_data_opD | 6'h4 ==
    decoder_inst_data_opD)); // @[Mux.scala 81:58]
  wire [32:0] decoder_inst_data_lo = {_decoder_inst_data_T_45,io_port_rdata}; // @[Cat.scala 31:58]
  wire [6:0] decoder_inst_data_hi = {_decoder_inst_data_T_17,_decoder_inst_data_T_27}; // @[Cat.scala 31:58]
  wire [39:0] decoder_inst_data = {_decoder_inst_data_T_17,_decoder_inst_data_T_27,_decoder_inst_data_T_45,io_port_rdata
    }; // @[Cat.scala 31:58]
  wire  _GEN_4 = 7'h1 == stage1_sram_addr_reg[11:5] ? lru_1 : lru_0; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_5 = 7'h2 == stage1_sram_addr_reg[11:5] ? lru_2 : _GEN_4; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_6 = 7'h3 == stage1_sram_addr_reg[11:5] ? lru_3 : _GEN_5; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_7 = 7'h4 == stage1_sram_addr_reg[11:5] ? lru_4 : _GEN_6; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_8 = 7'h5 == stage1_sram_addr_reg[11:5] ? lru_5 : _GEN_7; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_9 = 7'h6 == stage1_sram_addr_reg[11:5] ? lru_6 : _GEN_8; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_10 = 7'h7 == stage1_sram_addr_reg[11:5] ? lru_7 : _GEN_9; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_11 = 7'h8 == stage1_sram_addr_reg[11:5] ? lru_8 : _GEN_10; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_12 = 7'h9 == stage1_sram_addr_reg[11:5] ? lru_9 : _GEN_11; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_13 = 7'ha == stage1_sram_addr_reg[11:5] ? lru_10 : _GEN_12; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_14 = 7'hb == stage1_sram_addr_reg[11:5] ? lru_11 : _GEN_13; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_15 = 7'hc == stage1_sram_addr_reg[11:5] ? lru_12 : _GEN_14; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_16 = 7'hd == stage1_sram_addr_reg[11:5] ? lru_13 : _GEN_15; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_17 = 7'he == stage1_sram_addr_reg[11:5] ? lru_14 : _GEN_16; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_18 = 7'hf == stage1_sram_addr_reg[11:5] ? lru_15 : _GEN_17; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_19 = 7'h10 == stage1_sram_addr_reg[11:5] ? lru_16 : _GEN_18; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_20 = 7'h11 == stage1_sram_addr_reg[11:5] ? lru_17 : _GEN_19; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_21 = 7'h12 == stage1_sram_addr_reg[11:5] ? lru_18 : _GEN_20; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_22 = 7'h13 == stage1_sram_addr_reg[11:5] ? lru_19 : _GEN_21; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_23 = 7'h14 == stage1_sram_addr_reg[11:5] ? lru_20 : _GEN_22; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_24 = 7'h15 == stage1_sram_addr_reg[11:5] ? lru_21 : _GEN_23; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_25 = 7'h16 == stage1_sram_addr_reg[11:5] ? lru_22 : _GEN_24; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_26 = 7'h17 == stage1_sram_addr_reg[11:5] ? lru_23 : _GEN_25; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_27 = 7'h18 == stage1_sram_addr_reg[11:5] ? lru_24 : _GEN_26; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_28 = 7'h19 == stage1_sram_addr_reg[11:5] ? lru_25 : _GEN_27; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_29 = 7'h1a == stage1_sram_addr_reg[11:5] ? lru_26 : _GEN_28; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_30 = 7'h1b == stage1_sram_addr_reg[11:5] ? lru_27 : _GEN_29; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_31 = 7'h1c == stage1_sram_addr_reg[11:5] ? lru_28 : _GEN_30; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_32 = 7'h1d == stage1_sram_addr_reg[11:5] ? lru_29 : _GEN_31; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_33 = 7'h1e == stage1_sram_addr_reg[11:5] ? lru_30 : _GEN_32; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_34 = 7'h1f == stage1_sram_addr_reg[11:5] ? lru_31 : _GEN_33; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_35 = 7'h20 == stage1_sram_addr_reg[11:5] ? lru_32 : _GEN_34; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_36 = 7'h21 == stage1_sram_addr_reg[11:5] ? lru_33 : _GEN_35; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_37 = 7'h22 == stage1_sram_addr_reg[11:5] ? lru_34 : _GEN_36; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_38 = 7'h23 == stage1_sram_addr_reg[11:5] ? lru_35 : _GEN_37; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_39 = 7'h24 == stage1_sram_addr_reg[11:5] ? lru_36 : _GEN_38; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_40 = 7'h25 == stage1_sram_addr_reg[11:5] ? lru_37 : _GEN_39; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_41 = 7'h26 == stage1_sram_addr_reg[11:5] ? lru_38 : _GEN_40; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_42 = 7'h27 == stage1_sram_addr_reg[11:5] ? lru_39 : _GEN_41; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_43 = 7'h28 == stage1_sram_addr_reg[11:5] ? lru_40 : _GEN_42; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_44 = 7'h29 == stage1_sram_addr_reg[11:5] ? lru_41 : _GEN_43; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_45 = 7'h2a == stage1_sram_addr_reg[11:5] ? lru_42 : _GEN_44; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_46 = 7'h2b == stage1_sram_addr_reg[11:5] ? lru_43 : _GEN_45; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_47 = 7'h2c == stage1_sram_addr_reg[11:5] ? lru_44 : _GEN_46; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_48 = 7'h2d == stage1_sram_addr_reg[11:5] ? lru_45 : _GEN_47; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_49 = 7'h2e == stage1_sram_addr_reg[11:5] ? lru_46 : _GEN_48; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_50 = 7'h2f == stage1_sram_addr_reg[11:5] ? lru_47 : _GEN_49; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_51 = 7'h30 == stage1_sram_addr_reg[11:5] ? lru_48 : _GEN_50; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_52 = 7'h31 == stage1_sram_addr_reg[11:5] ? lru_49 : _GEN_51; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_53 = 7'h32 == stage1_sram_addr_reg[11:5] ? lru_50 : _GEN_52; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_54 = 7'h33 == stage1_sram_addr_reg[11:5] ? lru_51 : _GEN_53; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_55 = 7'h34 == stage1_sram_addr_reg[11:5] ? lru_52 : _GEN_54; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_56 = 7'h35 == stage1_sram_addr_reg[11:5] ? lru_53 : _GEN_55; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_57 = 7'h36 == stage1_sram_addr_reg[11:5] ? lru_54 : _GEN_56; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_58 = 7'h37 == stage1_sram_addr_reg[11:5] ? lru_55 : _GEN_57; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_59 = 7'h38 == stage1_sram_addr_reg[11:5] ? lru_56 : _GEN_58; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_60 = 7'h39 == stage1_sram_addr_reg[11:5] ? lru_57 : _GEN_59; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_61 = 7'h3a == stage1_sram_addr_reg[11:5] ? lru_58 : _GEN_60; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_62 = 7'h3b == stage1_sram_addr_reg[11:5] ? lru_59 : _GEN_61; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_63 = 7'h3c == stage1_sram_addr_reg[11:5] ? lru_60 : _GEN_62; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_64 = 7'h3d == stage1_sram_addr_reg[11:5] ? lru_61 : _GEN_63; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_65 = 7'h3e == stage1_sram_addr_reg[11:5] ? lru_62 : _GEN_64; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_66 = 7'h3f == stage1_sram_addr_reg[11:5] ? lru_63 : _GEN_65; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_67 = 7'h40 == stage1_sram_addr_reg[11:5] ? lru_64 : _GEN_66; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_68 = 7'h41 == stage1_sram_addr_reg[11:5] ? lru_65 : _GEN_67; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_69 = 7'h42 == stage1_sram_addr_reg[11:5] ? lru_66 : _GEN_68; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_70 = 7'h43 == stage1_sram_addr_reg[11:5] ? lru_67 : _GEN_69; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_71 = 7'h44 == stage1_sram_addr_reg[11:5] ? lru_68 : _GEN_70; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_72 = 7'h45 == stage1_sram_addr_reg[11:5] ? lru_69 : _GEN_71; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_73 = 7'h46 == stage1_sram_addr_reg[11:5] ? lru_70 : _GEN_72; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_74 = 7'h47 == stage1_sram_addr_reg[11:5] ? lru_71 : _GEN_73; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_75 = 7'h48 == stage1_sram_addr_reg[11:5] ? lru_72 : _GEN_74; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_76 = 7'h49 == stage1_sram_addr_reg[11:5] ? lru_73 : _GEN_75; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_77 = 7'h4a == stage1_sram_addr_reg[11:5] ? lru_74 : _GEN_76; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_78 = 7'h4b == stage1_sram_addr_reg[11:5] ? lru_75 : _GEN_77; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_79 = 7'h4c == stage1_sram_addr_reg[11:5] ? lru_76 : _GEN_78; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_80 = 7'h4d == stage1_sram_addr_reg[11:5] ? lru_77 : _GEN_79; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_81 = 7'h4e == stage1_sram_addr_reg[11:5] ? lru_78 : _GEN_80; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_82 = 7'h4f == stage1_sram_addr_reg[11:5] ? lru_79 : _GEN_81; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_83 = 7'h50 == stage1_sram_addr_reg[11:5] ? lru_80 : _GEN_82; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_84 = 7'h51 == stage1_sram_addr_reg[11:5] ? lru_81 : _GEN_83; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_85 = 7'h52 == stage1_sram_addr_reg[11:5] ? lru_82 : _GEN_84; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_86 = 7'h53 == stage1_sram_addr_reg[11:5] ? lru_83 : _GEN_85; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_87 = 7'h54 == stage1_sram_addr_reg[11:5] ? lru_84 : _GEN_86; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_88 = 7'h55 == stage1_sram_addr_reg[11:5] ? lru_85 : _GEN_87; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_89 = 7'h56 == stage1_sram_addr_reg[11:5] ? lru_86 : _GEN_88; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_90 = 7'h57 == stage1_sram_addr_reg[11:5] ? lru_87 : _GEN_89; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_91 = 7'h58 == stage1_sram_addr_reg[11:5] ? lru_88 : _GEN_90; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_92 = 7'h59 == stage1_sram_addr_reg[11:5] ? lru_89 : _GEN_91; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_93 = 7'h5a == stage1_sram_addr_reg[11:5] ? lru_90 : _GEN_92; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_94 = 7'h5b == stage1_sram_addr_reg[11:5] ? lru_91 : _GEN_93; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_95 = 7'h5c == stage1_sram_addr_reg[11:5] ? lru_92 : _GEN_94; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_96 = 7'h5d == stage1_sram_addr_reg[11:5] ? lru_93 : _GEN_95; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_97 = 7'h5e == stage1_sram_addr_reg[11:5] ? lru_94 : _GEN_96; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_98 = 7'h5f == stage1_sram_addr_reg[11:5] ? lru_95 : _GEN_97; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_99 = 7'h60 == stage1_sram_addr_reg[11:5] ? lru_96 : _GEN_98; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_100 = 7'h61 == stage1_sram_addr_reg[11:5] ? lru_97 : _GEN_99; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_101 = 7'h62 == stage1_sram_addr_reg[11:5] ? lru_98 : _GEN_100; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_102 = 7'h63 == stage1_sram_addr_reg[11:5] ? lru_99 : _GEN_101; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_103 = 7'h64 == stage1_sram_addr_reg[11:5] ? lru_100 : _GEN_102; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_104 = 7'h65 == stage1_sram_addr_reg[11:5] ? lru_101 : _GEN_103; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_105 = 7'h66 == stage1_sram_addr_reg[11:5] ? lru_102 : _GEN_104; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_106 = 7'h67 == stage1_sram_addr_reg[11:5] ? lru_103 : _GEN_105; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_107 = 7'h68 == stage1_sram_addr_reg[11:5] ? lru_104 : _GEN_106; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_108 = 7'h69 == stage1_sram_addr_reg[11:5] ? lru_105 : _GEN_107; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_109 = 7'h6a == stage1_sram_addr_reg[11:5] ? lru_106 : _GEN_108; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_110 = 7'h6b == stage1_sram_addr_reg[11:5] ? lru_107 : _GEN_109; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_111 = 7'h6c == stage1_sram_addr_reg[11:5] ? lru_108 : _GEN_110; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_112 = 7'h6d == stage1_sram_addr_reg[11:5] ? lru_109 : _GEN_111; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_113 = 7'h6e == stage1_sram_addr_reg[11:5] ? lru_110 : _GEN_112; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_114 = 7'h6f == stage1_sram_addr_reg[11:5] ? lru_111 : _GEN_113; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_115 = 7'h70 == stage1_sram_addr_reg[11:5] ? lru_112 : _GEN_114; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_116 = 7'h71 == stage1_sram_addr_reg[11:5] ? lru_113 : _GEN_115; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_117 = 7'h72 == stage1_sram_addr_reg[11:5] ? lru_114 : _GEN_116; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_118 = 7'h73 == stage1_sram_addr_reg[11:5] ? lru_115 : _GEN_117; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_119 = 7'h74 == stage1_sram_addr_reg[11:5] ? lru_116 : _GEN_118; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_120 = 7'h75 == stage1_sram_addr_reg[11:5] ? lru_117 : _GEN_119; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_121 = 7'h76 == stage1_sram_addr_reg[11:5] ? lru_118 : _GEN_120; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_122 = 7'h77 == stage1_sram_addr_reg[11:5] ? lru_119 : _GEN_121; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_123 = 7'h78 == stage1_sram_addr_reg[11:5] ? lru_120 : _GEN_122; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_124 = 7'h79 == stage1_sram_addr_reg[11:5] ? lru_121 : _GEN_123; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_125 = 7'h7a == stage1_sram_addr_reg[11:5] ? lru_122 : _GEN_124; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_126 = 7'h7b == stage1_sram_addr_reg[11:5] ? lru_123 : _GEN_125; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_127 = 7'h7c == stage1_sram_addr_reg[11:5] ? lru_124 : _GEN_126; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_128 = 7'h7d == stage1_sram_addr_reg[11:5] ? lru_125 : _GEN_127; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_129 = 7'h7e == stage1_sram_addr_reg[11:5] ? lru_126 : _GEN_128; // @[inst_cache.scala 187:{12,12}]
  wire  _GEN_130 = 7'h7f == stage1_sram_addr_reg[11:5] ? lru_127 : _GEN_129; // @[inst_cache.scala 187:{12,12}]
  wire  _lru_T_4 = _hit_T_3 ? 1'h0 : _GEN_130; // @[inst_cache.scala 187:12]
  wire  _lru_T_5 = _hit_T | _lru_T_4; // @[inst_cache.scala 186:12]
  wire  _lru_T_8 = ~_GEN_130; // @[inst_cache.scala 188:46]
  reg [31:0] stage2_sram_addr_reg; // @[inst_cache.scala 195:39]
  reg  stage2_sram_req_reg; // @[inst_cache.scala 205:38]
  reg  stage2_hit0_reg; // @[inst_cache.scala 209:34]
  reg [1:0] stage2_write_en_reg; // @[inst_cache.scala 227:38]
  wire  _stage2_write_en_reg_T_16 = access_stage1_sram_valid == 2'h1 ? 1'h0 : 1'h1; // @[inst_cache.scala 229:152]
  wire  _stage2_write_en_reg_T_17 = stage1_sram_req_reg ? _stage2_write_en_reg_T_16 : 1'h1; // @[inst_cache.scala 229:121]
  wire [39:0] icache_data_way0_0_rdata = icache_data_io_rdata; // @[inst_cache.scala 98:{36,36}]
  wire [39:0] icache_data_way0_1_rdata = icache_data_1_io_rdata; // @[inst_cache.scala 98:{36,36}]
  wire [39:0] _GEN_516 = 3'h1 == stage2_sram_addr_reg[4:2] ? icache_data_way0_1_rdata : icache_data_way0_0_rdata; // @[inst_cache.scala 238:{25,25}]
  wire [39:0] icache_data_way0_2_rdata = icache_data_2_io_rdata; // @[inst_cache.scala 98:{36,36}]
  wire [39:0] _GEN_517 = 3'h2 == stage2_sram_addr_reg[4:2] ? icache_data_way0_2_rdata : _GEN_516; // @[inst_cache.scala 238:{25,25}]
  wire [39:0] icache_data_way0_3_rdata = icache_data_3_io_rdata; // @[inst_cache.scala 98:{36,36}]
  wire [39:0] _GEN_518 = 3'h3 == stage2_sram_addr_reg[4:2] ? icache_data_way0_3_rdata : _GEN_517; // @[inst_cache.scala 238:{25,25}]
  wire [39:0] icache_data_way0_4_rdata = icache_data_4_io_rdata; // @[inst_cache.scala 98:{36,36}]
  wire [39:0] _GEN_519 = 3'h4 == stage2_sram_addr_reg[4:2] ? icache_data_way0_4_rdata : _GEN_518; // @[inst_cache.scala 238:{25,25}]
  wire [39:0] icache_data_way0_5_rdata = icache_data_5_io_rdata; // @[inst_cache.scala 98:{36,36}]
  wire [39:0] _GEN_520 = 3'h5 == stage2_sram_addr_reg[4:2] ? icache_data_way0_5_rdata : _GEN_519; // @[inst_cache.scala 238:{25,25}]
  wire [39:0] icache_data_way0_6_rdata = icache_data_6_io_rdata; // @[inst_cache.scala 98:{36,36}]
  wire [39:0] _GEN_521 = 3'h6 == stage2_sram_addr_reg[4:2] ? icache_data_way0_6_rdata : _GEN_520; // @[inst_cache.scala 238:{25,25}]
  wire [39:0] icache_data_way0_7_rdata = icache_data_7_io_rdata; // @[inst_cache.scala 98:{36,36}]
  wire [39:0] _GEN_522 = 3'h7 == stage2_sram_addr_reg[4:2] ? icache_data_way0_7_rdata : _GEN_521; // @[inst_cache.scala 238:{25,25}]
  wire [39:0] icache_data_way1_0_rdata = icache_data_8_io_rdata; // @[inst_cache.scala 99:{36,36}]
  wire [39:0] icache_data_way1_1_rdata = icache_data_9_io_rdata; // @[inst_cache.scala 99:{36,36}]
  wire [39:0] _GEN_524 = 3'h1 == stage2_sram_addr_reg[4:2] ? icache_data_way1_1_rdata : icache_data_way1_0_rdata; // @[inst_cache.scala 238:{25,25}]
  wire [39:0] icache_data_way1_2_rdata = icache_data_10_io_rdata; // @[inst_cache.scala 99:{36,36}]
  wire [39:0] _GEN_525 = 3'h2 == stage2_sram_addr_reg[4:2] ? icache_data_way1_2_rdata : _GEN_524; // @[inst_cache.scala 238:{25,25}]
  wire [39:0] icache_data_way1_3_rdata = icache_data_11_io_rdata; // @[inst_cache.scala 99:{36,36}]
  wire [39:0] _GEN_526 = 3'h3 == stage2_sram_addr_reg[4:2] ? icache_data_way1_3_rdata : _GEN_525; // @[inst_cache.scala 238:{25,25}]
  wire [39:0] icache_data_way1_4_rdata = icache_data_12_io_rdata; // @[inst_cache.scala 99:{36,36}]
  wire [39:0] _GEN_527 = 3'h4 == stage2_sram_addr_reg[4:2] ? icache_data_way1_4_rdata : _GEN_526; // @[inst_cache.scala 238:{25,25}]
  wire [39:0] icache_data_way1_5_rdata = icache_data_13_io_rdata; // @[inst_cache.scala 99:{36,36}]
  wire [39:0] _GEN_528 = 3'h5 == stage2_sram_addr_reg[4:2] ? icache_data_way1_5_rdata : _GEN_527; // @[inst_cache.scala 238:{25,25}]
  wire [39:0] icache_data_way1_6_rdata = icache_data_14_io_rdata; // @[inst_cache.scala 99:{36,36}]
  wire [39:0] _GEN_529 = 3'h6 == stage2_sram_addr_reg[4:2] ? icache_data_way1_6_rdata : _GEN_528; // @[inst_cache.scala 238:{25,25}]
  wire [39:0] icache_data_way1_7_rdata = icache_data_15_io_rdata; // @[inst_cache.scala 99:{36,36}]
  wire [39:0] _GEN_530 = 3'h7 == stage2_sram_addr_reg[4:2] ? icache_data_way1_7_rdata : _GEN_529; // @[inst_cache.scala 238:{25,25}]
  wire [39:0] hit_word_L = stage2_hit0_reg ? _GEN_522 : _GEN_530; // @[inst_cache.scala 238:25]
  reg  has_stage2_stall; // @[inst_cache.scala 240:35]
  reg [39:0] sram_rdata_L_Reg; // @[inst_cache.scala 243:35]
  wire [39:0] _access_sram_rdata_L_T_2 = _access_work_state_T_23 ? hit_word_L : 40'h0; // @[inst_cache.scala 246:84]
  wire [39:0] access_sram_rdata_L = _access_work_state_T_8 ? wait_data_L : _access_sram_rdata_L_T_2; // @[inst_cache.scala 246:35]
  wire  _wait_data_L_T_3 = write_counter == 3'h0; // @[inst_cache.scala 278:100]
  wire  _wait_data_L_T_7 = _access_work_state_T_38 & io_port_rvalid; // @[inst_cache.scala 279:53]
  wire [2:0] _write_counter_T_8 = write_counter + 3'h1; // @[inst_cache.scala 284:195]
  wire  _icache_data_way0_0_wen_T_7 = _wait_data_L_T_7 & _lru_T_8 & _wait_data_L_T_3; // @[inst_cache.scala 291:52]
  wire  _icache_data_way0_1_wen_T_6 = write_counter == 3'h1; // @[inst_cache.scala 291:69]
  wire  _icache_data_way0_1_wen_T_7 = _wait_data_L_T_7 & _lru_T_8 & write_counter == 3'h1; // @[inst_cache.scala 291:52]
  wire  _icache_data_way0_2_wen_T_6 = write_counter == 3'h2; // @[inst_cache.scala 291:69]
  wire  _icache_data_way0_2_wen_T_7 = _wait_data_L_T_7 & _lru_T_8 & write_counter == 3'h2; // @[inst_cache.scala 291:52]
  wire  _icache_data_way0_3_wen_T_6 = write_counter == 3'h3; // @[inst_cache.scala 291:69]
  wire  _icache_data_way0_3_wen_T_7 = _wait_data_L_T_7 & _lru_T_8 & write_counter == 3'h3; // @[inst_cache.scala 291:52]
  wire  _icache_data_way0_4_wen_T_6 = write_counter == 3'h4; // @[inst_cache.scala 291:69]
  wire  _icache_data_way0_4_wen_T_7 = _wait_data_L_T_7 & _lru_T_8 & write_counter == 3'h4; // @[inst_cache.scala 291:52]
  wire  _icache_data_way0_5_wen_T_6 = write_counter == 3'h5; // @[inst_cache.scala 291:69]
  wire  _icache_data_way0_5_wen_T_7 = _wait_data_L_T_7 & _lru_T_8 & write_counter == 3'h5; // @[inst_cache.scala 291:52]
  wire  _icache_data_way0_6_wen_T_6 = write_counter == 3'h6; // @[inst_cache.scala 291:69]
  wire  _icache_data_way0_6_wen_T_7 = _wait_data_L_T_7 & _lru_T_8 & write_counter == 3'h6; // @[inst_cache.scala 291:52]
  wire  _icache_data_way0_7_wen_T_6 = write_counter == 3'h7; // @[inst_cache.scala 291:69]
  wire  _icache_data_way0_7_wen_T_7 = _wait_data_L_T_7 & _lru_T_8 & write_counter == 3'h7; // @[inst_cache.scala 291:52]
  wire  _icache_data_way1_0_wen_T_7 = _wait_data_L_T_7 & _GEN_130 & _wait_data_L_T_3; // @[inst_cache.scala 293:52]
  wire  _icache_data_way1_1_wen_T_7 = _wait_data_L_T_7 & _GEN_130 & _icache_data_way0_1_wen_T_6; // @[inst_cache.scala 293:52]
  wire  _icache_data_way1_2_wen_T_7 = _wait_data_L_T_7 & _GEN_130 & _icache_data_way0_2_wen_T_6; // @[inst_cache.scala 293:52]
  wire  _icache_data_way1_3_wen_T_7 = _wait_data_L_T_7 & _GEN_130 & _icache_data_way0_3_wen_T_6; // @[inst_cache.scala 293:52]
  wire  _icache_data_way1_4_wen_T_7 = _wait_data_L_T_7 & _GEN_130 & _icache_data_way0_4_wen_T_6; // @[inst_cache.scala 293:52]
  wire  _icache_data_way1_5_wen_T_7 = _wait_data_L_T_7 & _GEN_130 & _icache_data_way0_5_wen_T_6; // @[inst_cache.scala 293:52]
  wire  _icache_data_way1_6_wen_T_7 = _wait_data_L_T_7 & _GEN_130 & _icache_data_way0_6_wen_T_6; // @[inst_cache.scala 293:52]
  wire  _icache_data_way1_7_wen_T_7 = _wait_data_L_T_7 & _GEN_130 & _icache_data_way0_7_wen_T_6; // @[inst_cache.scala 293:52]
  wire [20:0] _T_13 = {1'h1,stage1_sram_addr_reg[31:12]}; // @[Cat.scala 31:58]
  wire [31:0] _io_port_araddr_T_3 = {stage1_sram_phy_addr_reg[31:5],5'h0}; // @[Cat.scala 31:58]
  wire [31:0] _io_port_araddr_T_4 = _access_work_state_T_35 ? _io_port_araddr_T_3 : 32'h0; // @[inst_cache.scala 308:12]
  wire [2:0] _io_port_arlen_T_1 = stage1_sram_cache_reg ? 3'h7 : 3'h0; // @[inst_cache.scala 310:26]
  wire  _io_port_sram_write_en_T_3 = ~stage2_sram_req_reg & stage2_sram_addr_reg[1:0] != 2'h0; // @[inst_cache.scala 345:31]
  wire [1:0] _io_port_sram_write_en_T_5 = stage2_sram_req_reg | _io_port_sram_write_en_T_3 ? stage2_write_en_reg : 2'h0; // @[inst_cache.scala 344:62]
  icache_tag icache_tag ( // @[inst_cache.scala 93:34]
    .clock(icache_tag_clock),
    .reset(icache_tag_reset),
    .io_wen(icache_tag_io_wen),
    .io_wdata(icache_tag_io_wdata),
    .io_addr(icache_tag_io_addr),
    .io_hit(icache_tag_io_hit),
    .io_valid(icache_tag_io_valid),
    .io_asid(icache_tag_io_asid)
  );
  icache_tag icache_tag_1 ( // @[inst_cache.scala 95:34]
    .clock(icache_tag_1_clock),
    .reset(icache_tag_1_reset),
    .io_wen(icache_tag_1_io_wen),
    .io_wdata(icache_tag_1_io_wdata),
    .io_addr(icache_tag_1_io_addr),
    .io_hit(icache_tag_1_io_hit),
    .io_valid(icache_tag_1_io_valid),
    .io_asid(icache_tag_1_io_asid)
  );
  icache_data icache_data ( // @[inst_cache.scala 98:55]
    .clock(icache_data_clock),
    .io_wen(icache_data_io_wen),
    .io_addr(icache_data_io_addr),
    .io_wdata(icache_data_io_wdata),
    .io_rdata(icache_data_io_rdata)
  );
  icache_data icache_data_1 ( // @[inst_cache.scala 98:55]
    .clock(icache_data_1_clock),
    .io_wen(icache_data_1_io_wen),
    .io_addr(icache_data_1_io_addr),
    .io_wdata(icache_data_1_io_wdata),
    .io_rdata(icache_data_1_io_rdata)
  );
  icache_data icache_data_2 ( // @[inst_cache.scala 98:55]
    .clock(icache_data_2_clock),
    .io_wen(icache_data_2_io_wen),
    .io_addr(icache_data_2_io_addr),
    .io_wdata(icache_data_2_io_wdata),
    .io_rdata(icache_data_2_io_rdata)
  );
  icache_data icache_data_3 ( // @[inst_cache.scala 98:55]
    .clock(icache_data_3_clock),
    .io_wen(icache_data_3_io_wen),
    .io_addr(icache_data_3_io_addr),
    .io_wdata(icache_data_3_io_wdata),
    .io_rdata(icache_data_3_io_rdata)
  );
  icache_data icache_data_4 ( // @[inst_cache.scala 98:55]
    .clock(icache_data_4_clock),
    .io_wen(icache_data_4_io_wen),
    .io_addr(icache_data_4_io_addr),
    .io_wdata(icache_data_4_io_wdata),
    .io_rdata(icache_data_4_io_rdata)
  );
  icache_data icache_data_5 ( // @[inst_cache.scala 98:55]
    .clock(icache_data_5_clock),
    .io_wen(icache_data_5_io_wen),
    .io_addr(icache_data_5_io_addr),
    .io_wdata(icache_data_5_io_wdata),
    .io_rdata(icache_data_5_io_rdata)
  );
  icache_data icache_data_6 ( // @[inst_cache.scala 98:55]
    .clock(icache_data_6_clock),
    .io_wen(icache_data_6_io_wen),
    .io_addr(icache_data_6_io_addr),
    .io_wdata(icache_data_6_io_wdata),
    .io_rdata(icache_data_6_io_rdata)
  );
  icache_data icache_data_7 ( // @[inst_cache.scala 98:55]
    .clock(icache_data_7_clock),
    .io_wen(icache_data_7_io_wen),
    .io_addr(icache_data_7_io_addr),
    .io_wdata(icache_data_7_io_wdata),
    .io_rdata(icache_data_7_io_rdata)
  );
  icache_data icache_data_8 ( // @[inst_cache.scala 99:55]
    .clock(icache_data_8_clock),
    .io_wen(icache_data_8_io_wen),
    .io_addr(icache_data_8_io_addr),
    .io_wdata(icache_data_8_io_wdata),
    .io_rdata(icache_data_8_io_rdata)
  );
  icache_data icache_data_9 ( // @[inst_cache.scala 99:55]
    .clock(icache_data_9_clock),
    .io_wen(icache_data_9_io_wen),
    .io_addr(icache_data_9_io_addr),
    .io_wdata(icache_data_9_io_wdata),
    .io_rdata(icache_data_9_io_rdata)
  );
  icache_data icache_data_10 ( // @[inst_cache.scala 99:55]
    .clock(icache_data_10_clock),
    .io_wen(icache_data_10_io_wen),
    .io_addr(icache_data_10_io_addr),
    .io_wdata(icache_data_10_io_wdata),
    .io_rdata(icache_data_10_io_rdata)
  );
  icache_data icache_data_11 ( // @[inst_cache.scala 99:55]
    .clock(icache_data_11_clock),
    .io_wen(icache_data_11_io_wen),
    .io_addr(icache_data_11_io_addr),
    .io_wdata(icache_data_11_io_wdata),
    .io_rdata(icache_data_11_io_rdata)
  );
  icache_data icache_data_12 ( // @[inst_cache.scala 99:55]
    .clock(icache_data_12_clock),
    .io_wen(icache_data_12_io_wen),
    .io_addr(icache_data_12_io_addr),
    .io_wdata(icache_data_12_io_wdata),
    .io_rdata(icache_data_12_io_rdata)
  );
  icache_data icache_data_13 ( // @[inst_cache.scala 99:55]
    .clock(icache_data_13_clock),
    .io_wen(icache_data_13_io_wen),
    .io_addr(icache_data_13_io_addr),
    .io_wdata(icache_data_13_io_wdata),
    .io_rdata(icache_data_13_io_rdata)
  );
  icache_data icache_data_14 ( // @[inst_cache.scala 99:55]
    .clock(icache_data_14_clock),
    .io_wen(icache_data_14_io_wen),
    .io_addr(icache_data_14_io_addr),
    .io_wdata(icache_data_14_io_wdata),
    .io_rdata(icache_data_14_io_rdata)
  );
  icache_data icache_data_15 ( // @[inst_cache.scala 99:55]
    .clock(icache_data_15_clock),
    .io_wen(icache_data_15_io_wen),
    .io_addr(icache_data_15_io_addr),
    .io_wdata(icache_data_15_io_wdata),
    .io_rdata(icache_data_15_io_rdata)
  );
  assign io_port_araddr = _access_work_state_T ? stage1_sram_phy_addr_reg : _io_port_araddr_T_4; // @[inst_cache.scala 307:26]
  assign io_port_arlen = {{1'd0}, _io_port_arlen_T_1}; // @[inst_cache.scala 310:20]
  assign io_port_arburst = {{1'd0}, stage1_sram_cache_reg}; // @[inst_cache.scala 312:21]
  assign io_port_arvalid = (_access_work_state_T | _access_work_state_T_35) & stage1_exception == 2'h0; // @[inst_cache.scala 317:102]
  assign io_port_sram_write_en = io_inst_buffer_full ? 2'h0 : _io_port_sram_write_en_T_5; // @[inst_cache.scala 344:33]
  assign io_port_sram_rdata_L = _stage2_stall_T_5 & has_stage2_stall ? access_sram_rdata_L : sram_rdata_L_Reg; // @[inst_cache.scala 253:32]
  assign io_stage2_stall = (access_work_state == 4'h1 | access_work_state == 4'h4 | stage1_exception != 2'h0) &
    _stage2_stall_T_5; // @[inst_cache.scala 156:129]
  assign io_stage2_exception = stage2_exception; // @[inst_cache.scala 304:25]
  assign io_v_addr_for_tlb = stage1_sram_addr_reg; // @[inst_cache.scala 145:23]
  assign io_tlb_req = ~stage1_sram_addr_reg[31] | stage1_sram_addr_reg[31:30] == 2'h3; // @[macros.scala 424:18]
  assign icache_tag_clock = clock;
  assign icache_tag_reset = reset;
  assign icache_tag_io_wen = _stage1_finished_T_1 & _lru_T_8; // @[inst_cache.scala 295:62]
  assign icache_tag_io_wdata = _stage1_finished_T_1 ? _T_13 : 21'h0; // @[inst_cache.scala 297:30]
  assign icache_tag_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 166:25]
  assign icache_tag_io_asid = io_cp0_asid; // @[inst_cache.scala 94:23]
  assign icache_tag_1_clock = clock;
  assign icache_tag_1_reset = reset;
  assign icache_tag_1_io_wen = _stage1_finished_T_1 & _GEN_130; // @[inst_cache.scala 296:63]
  assign icache_tag_1_io_wdata = _stage1_finished_T_1 ? _T_13 : 21'h0; // @[inst_cache.scala 298:30]
  assign icache_tag_1_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 167:25]
  assign icache_tag_1_io_asid = io_cp0_asid; // @[inst_cache.scala 96:23]
  assign icache_data_clock = clock;
  assign icache_data_io_wen = _icache_data_way0_0_wen_T_7 ? 5'h1f : 5'h0; // @[inst_cache.scala 290:55]
  assign icache_data_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 172:34 98:36]
  assign icache_data_io_wdata = {decoder_inst_data_hi,decoder_inst_data_lo}; // @[Cat.scala 31:58]
  assign icache_data_1_clock = clock;
  assign icache_data_1_io_wen = _icache_data_way0_1_wen_T_7 ? 5'h1f : 5'h0; // @[inst_cache.scala 290:55]
  assign icache_data_1_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 172:34 98:36]
  assign icache_data_1_io_wdata = {decoder_inst_data_hi,decoder_inst_data_lo}; // @[Cat.scala 31:58]
  assign icache_data_2_clock = clock;
  assign icache_data_2_io_wen = _icache_data_way0_2_wen_T_7 ? 5'h1f : 5'h0; // @[inst_cache.scala 290:55]
  assign icache_data_2_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 172:34 98:36]
  assign icache_data_2_io_wdata = {decoder_inst_data_hi,decoder_inst_data_lo}; // @[Cat.scala 31:58]
  assign icache_data_3_clock = clock;
  assign icache_data_3_io_wen = _icache_data_way0_3_wen_T_7 ? 5'h1f : 5'h0; // @[inst_cache.scala 290:55]
  assign icache_data_3_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 172:34 98:36]
  assign icache_data_3_io_wdata = {decoder_inst_data_hi,decoder_inst_data_lo}; // @[Cat.scala 31:58]
  assign icache_data_4_clock = clock;
  assign icache_data_4_io_wen = _icache_data_way0_4_wen_T_7 ? 5'h1f : 5'h0; // @[inst_cache.scala 290:55]
  assign icache_data_4_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 172:34 98:36]
  assign icache_data_4_io_wdata = {decoder_inst_data_hi,decoder_inst_data_lo}; // @[Cat.scala 31:58]
  assign icache_data_5_clock = clock;
  assign icache_data_5_io_wen = _icache_data_way0_5_wen_T_7 ? 5'h1f : 5'h0; // @[inst_cache.scala 290:55]
  assign icache_data_5_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 172:34 98:36]
  assign icache_data_5_io_wdata = {decoder_inst_data_hi,decoder_inst_data_lo}; // @[Cat.scala 31:58]
  assign icache_data_6_clock = clock;
  assign icache_data_6_io_wen = _icache_data_way0_6_wen_T_7 ? 5'h1f : 5'h0; // @[inst_cache.scala 290:55]
  assign icache_data_6_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 172:34 98:36]
  assign icache_data_6_io_wdata = {decoder_inst_data_hi,decoder_inst_data_lo}; // @[Cat.scala 31:58]
  assign icache_data_7_clock = clock;
  assign icache_data_7_io_wen = _icache_data_way0_7_wen_T_7 ? 5'h1f : 5'h0; // @[inst_cache.scala 290:55]
  assign icache_data_7_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 172:34 98:36]
  assign icache_data_7_io_wdata = {decoder_inst_data_hi,decoder_inst_data_lo}; // @[Cat.scala 31:58]
  assign icache_data_8_clock = clock;
  assign icache_data_8_io_wen = _icache_data_way1_0_wen_T_7 ? 5'h1f : 5'h0; // @[inst_cache.scala 292:55]
  assign icache_data_8_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 177:34 99:36]
  assign icache_data_8_io_wdata = {decoder_inst_data_hi,decoder_inst_data_lo}; // @[Cat.scala 31:58]
  assign icache_data_9_clock = clock;
  assign icache_data_9_io_wen = _icache_data_way1_1_wen_T_7 ? 5'h1f : 5'h0; // @[inst_cache.scala 292:55]
  assign icache_data_9_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 177:34 99:36]
  assign icache_data_9_io_wdata = {decoder_inst_data_hi,decoder_inst_data_lo}; // @[Cat.scala 31:58]
  assign icache_data_10_clock = clock;
  assign icache_data_10_io_wen = _icache_data_way1_2_wen_T_7 ? 5'h1f : 5'h0; // @[inst_cache.scala 292:55]
  assign icache_data_10_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 177:34 99:36]
  assign icache_data_10_io_wdata = {decoder_inst_data_hi,decoder_inst_data_lo}; // @[Cat.scala 31:58]
  assign icache_data_11_clock = clock;
  assign icache_data_11_io_wen = _icache_data_way1_3_wen_T_7 ? 5'h1f : 5'h0; // @[inst_cache.scala 292:55]
  assign icache_data_11_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 177:34 99:36]
  assign icache_data_11_io_wdata = {decoder_inst_data_hi,decoder_inst_data_lo}; // @[Cat.scala 31:58]
  assign icache_data_12_clock = clock;
  assign icache_data_12_io_wen = _icache_data_way1_4_wen_T_7 ? 5'h1f : 5'h0; // @[inst_cache.scala 292:55]
  assign icache_data_12_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 177:34 99:36]
  assign icache_data_12_io_wdata = {decoder_inst_data_hi,decoder_inst_data_lo}; // @[Cat.scala 31:58]
  assign icache_data_13_clock = clock;
  assign icache_data_13_io_wen = _icache_data_way1_5_wen_T_7 ? 5'h1f : 5'h0; // @[inst_cache.scala 292:55]
  assign icache_data_13_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 177:34 99:36]
  assign icache_data_13_io_wdata = {decoder_inst_data_hi,decoder_inst_data_lo}; // @[Cat.scala 31:58]
  assign icache_data_14_clock = clock;
  assign icache_data_14_io_wen = _icache_data_way1_6_wen_T_7 ? 5'h1f : 5'h0; // @[inst_cache.scala 292:55]
  assign icache_data_14_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 177:34 99:36]
  assign icache_data_14_io_wdata = {decoder_inst_data_hi,decoder_inst_data_lo}; // @[Cat.scala 31:58]
  assign icache_data_15_clock = clock;
  assign icache_data_15_io_wen = _icache_data_way1_7_wen_T_7 ? 5'h1f : 5'h0; // @[inst_cache.scala 292:55]
  assign icache_data_15_io_addr = stage1_sram_addr_reg; // @[inst_cache.scala 177:34 99:36]
  assign icache_data_15_io_wdata = {decoder_inst_data_hi,decoder_inst_data_lo}; // @[Cat.scala 31:58]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_0 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h0 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_0 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_0 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_0 <= lru_127;
      end else begin
        lru_0 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_1 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h1 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_1 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_1 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_1 <= lru_127;
      end else begin
        lru_1 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_2 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h2 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_2 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_2 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_2 <= lru_127;
      end else begin
        lru_2 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_3 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h3 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_3 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_3 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_3 <= lru_127;
      end else begin
        lru_3 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_4 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h4 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_4 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_4 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_4 <= lru_127;
      end else begin
        lru_4 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_5 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h5 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_5 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_5 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_5 <= lru_127;
      end else begin
        lru_5 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_6 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h6 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_6 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_6 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_6 <= lru_127;
      end else begin
        lru_6 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_7 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h7 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_7 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_7 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_7 <= lru_127;
      end else begin
        lru_7 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_8 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h8 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_8 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_8 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_8 <= lru_127;
      end else begin
        lru_8 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_9 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h9 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_9 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_9 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_9 <= lru_127;
      end else begin
        lru_9 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_10 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'ha == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_10 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_10 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_10 <= lru_127;
      end else begin
        lru_10 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_11 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'hb == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_11 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_11 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_11 <= lru_127;
      end else begin
        lru_11 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_12 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'hc == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_12 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_12 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_12 <= lru_127;
      end else begin
        lru_12 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_13 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'hd == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_13 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_13 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_13 <= lru_127;
      end else begin
        lru_13 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_14 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'he == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_14 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_14 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_14 <= lru_127;
      end else begin
        lru_14 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_15 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'hf == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_15 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_15 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_15 <= lru_127;
      end else begin
        lru_15 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_16 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h10 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_16 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_16 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_16 <= lru_127;
      end else begin
        lru_16 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_17 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h11 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_17 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_17 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_17 <= lru_127;
      end else begin
        lru_17 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_18 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h12 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_18 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_18 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_18 <= lru_127;
      end else begin
        lru_18 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_19 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h13 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_19 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_19 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_19 <= lru_127;
      end else begin
        lru_19 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_20 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h14 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_20 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_20 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_20 <= lru_127;
      end else begin
        lru_20 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_21 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h15 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_21 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_21 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_21 <= lru_127;
      end else begin
        lru_21 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_22 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h16 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_22 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_22 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_22 <= lru_127;
      end else begin
        lru_22 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_23 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h17 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_23 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_23 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_23 <= lru_127;
      end else begin
        lru_23 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_24 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h18 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_24 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_24 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_24 <= lru_127;
      end else begin
        lru_24 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_25 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h19 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_25 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_25 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_25 <= lru_127;
      end else begin
        lru_25 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_26 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h1a == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_26 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_26 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_26 <= lru_127;
      end else begin
        lru_26 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_27 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h1b == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_27 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_27 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_27 <= lru_127;
      end else begin
        lru_27 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_28 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h1c == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_28 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_28 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_28 <= lru_127;
      end else begin
        lru_28 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_29 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h1d == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_29 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_29 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_29 <= lru_127;
      end else begin
        lru_29 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_30 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h1e == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_30 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_30 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_30 <= lru_127;
      end else begin
        lru_30 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_31 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h1f == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_31 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_31 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_31 <= lru_127;
      end else begin
        lru_31 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_32 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h20 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_32 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_32 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_32 <= lru_127;
      end else begin
        lru_32 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_33 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h21 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_33 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_33 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_33 <= lru_127;
      end else begin
        lru_33 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_34 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h22 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_34 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_34 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_34 <= lru_127;
      end else begin
        lru_34 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_35 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h23 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_35 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_35 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_35 <= lru_127;
      end else begin
        lru_35 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_36 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h24 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_36 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_36 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_36 <= lru_127;
      end else begin
        lru_36 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_37 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h25 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_37 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_37 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_37 <= lru_127;
      end else begin
        lru_37 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_38 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h26 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_38 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_38 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_38 <= lru_127;
      end else begin
        lru_38 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_39 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h27 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_39 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_39 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_39 <= lru_127;
      end else begin
        lru_39 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_40 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h28 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_40 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_40 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_40 <= lru_127;
      end else begin
        lru_40 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_41 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h29 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_41 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_41 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_41 <= lru_127;
      end else begin
        lru_41 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_42 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h2a == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_42 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_42 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_42 <= lru_127;
      end else begin
        lru_42 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_43 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h2b == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_43 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_43 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_43 <= lru_127;
      end else begin
        lru_43 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_44 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h2c == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_44 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_44 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_44 <= lru_127;
      end else begin
        lru_44 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_45 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h2d == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_45 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_45 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_45 <= lru_127;
      end else begin
        lru_45 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_46 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h2e == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_46 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_46 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_46 <= lru_127;
      end else begin
        lru_46 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_47 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h2f == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_47 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_47 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_47 <= lru_127;
      end else begin
        lru_47 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_48 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h30 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_48 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_48 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_48 <= lru_127;
      end else begin
        lru_48 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_49 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h31 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_49 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_49 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_49 <= lru_127;
      end else begin
        lru_49 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_50 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h32 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_50 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_50 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_50 <= lru_127;
      end else begin
        lru_50 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_51 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h33 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_51 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_51 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_51 <= lru_127;
      end else begin
        lru_51 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_52 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h34 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_52 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_52 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_52 <= lru_127;
      end else begin
        lru_52 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_53 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h35 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_53 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_53 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_53 <= lru_127;
      end else begin
        lru_53 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_54 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h36 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_54 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_54 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_54 <= lru_127;
      end else begin
        lru_54 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_55 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h37 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_55 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_55 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_55 <= lru_127;
      end else begin
        lru_55 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_56 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h38 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_56 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_56 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_56 <= lru_127;
      end else begin
        lru_56 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_57 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h39 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_57 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_57 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_57 <= lru_127;
      end else begin
        lru_57 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_58 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h3a == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_58 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_58 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_58 <= lru_127;
      end else begin
        lru_58 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_59 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h3b == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_59 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_59 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_59 <= lru_127;
      end else begin
        lru_59 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_60 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h3c == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_60 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_60 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_60 <= lru_127;
      end else begin
        lru_60 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_61 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h3d == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_61 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_61 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_61 <= lru_127;
      end else begin
        lru_61 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_62 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h3e == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_62 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_62 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_62 <= lru_127;
      end else begin
        lru_62 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_63 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h3f == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_63 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_63 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_63 <= lru_127;
      end else begin
        lru_63 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_64 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h40 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_64 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_64 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_64 <= lru_127;
      end else begin
        lru_64 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_65 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h41 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_65 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_65 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_65 <= lru_127;
      end else begin
        lru_65 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_66 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h42 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_66 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_66 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_66 <= lru_127;
      end else begin
        lru_66 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_67 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h43 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_67 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_67 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_67 <= lru_127;
      end else begin
        lru_67 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_68 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h44 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_68 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_68 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_68 <= lru_127;
      end else begin
        lru_68 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_69 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h45 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_69 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_69 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_69 <= lru_127;
      end else begin
        lru_69 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_70 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h46 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_70 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_70 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_70 <= lru_127;
      end else begin
        lru_70 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_71 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h47 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_71 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_71 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_71 <= lru_127;
      end else begin
        lru_71 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_72 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h48 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_72 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_72 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_72 <= lru_127;
      end else begin
        lru_72 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_73 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h49 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_73 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_73 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_73 <= lru_127;
      end else begin
        lru_73 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_74 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h4a == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_74 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_74 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_74 <= lru_127;
      end else begin
        lru_74 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_75 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h4b == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_75 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_75 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_75 <= lru_127;
      end else begin
        lru_75 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_76 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h4c == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_76 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_76 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_76 <= lru_127;
      end else begin
        lru_76 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_77 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h4d == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_77 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_77 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_77 <= lru_127;
      end else begin
        lru_77 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_78 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h4e == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_78 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_78 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_78 <= lru_127;
      end else begin
        lru_78 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_79 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h4f == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_79 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_79 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_79 <= lru_127;
      end else begin
        lru_79 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_80 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h50 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_80 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_80 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_80 <= lru_127;
      end else begin
        lru_80 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_81 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h51 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_81 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_81 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_81 <= lru_127;
      end else begin
        lru_81 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_82 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h52 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_82 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_82 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_82 <= lru_127;
      end else begin
        lru_82 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_83 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h53 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_83 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_83 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_83 <= lru_127;
      end else begin
        lru_83 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_84 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h54 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_84 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_84 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_84 <= lru_127;
      end else begin
        lru_84 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_85 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h55 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_85 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_85 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_85 <= lru_127;
      end else begin
        lru_85 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_86 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h56 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_86 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_86 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_86 <= lru_127;
      end else begin
        lru_86 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_87 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h57 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_87 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_87 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_87 <= lru_127;
      end else begin
        lru_87 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_88 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h58 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_88 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_88 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_88 <= lru_127;
      end else begin
        lru_88 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_89 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h59 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_89 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_89 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_89 <= lru_127;
      end else begin
        lru_89 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_90 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h5a == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_90 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_90 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_90 <= lru_127;
      end else begin
        lru_90 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_91 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h5b == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_91 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_91 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_91 <= lru_127;
      end else begin
        lru_91 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_92 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h5c == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_92 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_92 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_92 <= lru_127;
      end else begin
        lru_92 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_93 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h5d == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_93 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_93 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_93 <= lru_127;
      end else begin
        lru_93 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_94 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h5e == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_94 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_94 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_94 <= lru_127;
      end else begin
        lru_94 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_95 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h5f == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_95 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_95 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_95 <= lru_127;
      end else begin
        lru_95 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_96 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h60 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_96 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_96 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_96 <= lru_127;
      end else begin
        lru_96 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_97 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h61 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_97 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_97 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_97 <= lru_127;
      end else begin
        lru_97 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_98 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h62 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_98 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_98 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_98 <= lru_127;
      end else begin
        lru_98 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_99 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h63 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_99 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_99 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_99 <= lru_127;
      end else begin
        lru_99 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_100 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h64 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_100 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_100 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_100 <= lru_127;
      end else begin
        lru_100 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_101 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h65 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_101 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_101 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_101 <= lru_127;
      end else begin
        lru_101 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_102 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h66 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_102 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_102 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_102 <= lru_127;
      end else begin
        lru_102 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_103 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h67 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_103 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_103 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_103 <= lru_127;
      end else begin
        lru_103 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_104 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h68 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_104 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_104 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_104 <= lru_127;
      end else begin
        lru_104 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_105 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h69 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_105 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_105 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_105 <= lru_127;
      end else begin
        lru_105 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_106 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h6a == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_106 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_106 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_106 <= lru_127;
      end else begin
        lru_106 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_107 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h6b == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_107 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_107 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_107 <= lru_127;
      end else begin
        lru_107 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_108 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h6c == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_108 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_108 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_108 <= lru_127;
      end else begin
        lru_108 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_109 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h6d == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_109 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_109 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_109 <= lru_127;
      end else begin
        lru_109 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_110 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h6e == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_110 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_110 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_110 <= lru_127;
      end else begin
        lru_110 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_111 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h6f == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_111 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_111 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_111 <= lru_127;
      end else begin
        lru_111 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_112 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h70 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_112 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_112 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_112 <= lru_127;
      end else begin
        lru_112 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_113 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h71 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_113 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_113 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_113 <= lru_127;
      end else begin
        lru_113 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_114 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h72 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_114 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_114 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_114 <= lru_127;
      end else begin
        lru_114 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_115 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h73 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_115 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_115 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_115 <= lru_127;
      end else begin
        lru_115 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_116 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h74 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_116 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_116 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_116 <= lru_127;
      end else begin
        lru_116 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_117 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h75 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_117 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_117 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_117 <= lru_127;
      end else begin
        lru_117 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_118 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h76 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_118 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_118 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_118 <= lru_127;
      end else begin
        lru_118 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_119 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h77 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_119 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_119 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_119 <= lru_127;
      end else begin
        lru_119 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_120 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h78 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_120 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_120 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_120 <= lru_127;
      end else begin
        lru_120 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_121 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h79 == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_121 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_121 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_121 <= lru_127;
      end else begin
        lru_121 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_122 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h7a == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_122 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_122 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_122 <= lru_127;
      end else begin
        lru_122 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_123 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h7b == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_123 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_123 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_123 <= lru_127;
      end else begin
        lru_123 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_124 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h7c == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_124 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_124 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_124 <= lru_127;
      end else begin
        lru_124 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_125 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h7d == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_125 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_125 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_125 <= lru_127;
      end else begin
        lru_125 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_126 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h7e == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_126 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_126 <= ~_GEN_130;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_126 <= lru_127;
      end else begin
        lru_126 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 185:37]
      lru_127 <= 1'h0; // @[inst_cache.scala 185:43 187:{12,12} 188:12]
    end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin // @[inst_cache.scala 86:22]
      if (_stage2_stall_T) begin
        lru_127 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_127 <= ~_GEN_130;
      end else if (!(7'h7f == stage1_sram_addr_reg[11:5])) begin
        lru_127 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 276:22]
      work_state <= 4'h1;
    end else if (_stage2_stall_T_3) begin // @[inst_cache.scala 256:30]
      work_state <= 4'h1;
    end else if (work_state == 4'h2 & io_port_arready) begin // @[inst_cache.scala 257:12]
      work_state <= 4'h3;
    end else if (_stage1_finished_T_2) begin // @[inst_cache.scala 258:12]
      work_state <= {{1'd0}, _access_work_state_T_7};
    end else if (work_state == 4'h4) begin
      work_state <= {{1'd0}, _access_work_state_T_22};
    end else begin
      work_state <= _access_work_state_T_47;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 284:25]
      write_counter <= 3'h0; // @[inst_cache.scala 284:{105,159}]
    end else if (_access_work_state_T_38 | _stage1_finished_T_2) begin
      if (io_port_rvalid & io_port_rlast) begin
        write_counter <= 3'h0;
      end else if (io_port_rvalid) begin
        write_counter <= _write_counter_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 278:23]
      wait_data_L <= 40'h0;
    end else if (_stage1_finished_T_2 & io_port_rvalid & write_counter == 3'h0) begin // @[inst_cache.scala 279:13]
      wait_data_L <= decoder_inst_data;
    end else if (_access_work_state_T_38 & io_port_rvalid & write_counter == stage1_sram_addr_reg[4:2]) begin
      wait_data_L <= decoder_inst_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 121:18 89:28]
      stage1_stall_reg <= 1'h0;
    end else begin
      stage1_stall_reg <= io_port_sram_req;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      stage1_sram_addr_reg <= 32'h0; // @[Reg.scala 29:22]
    end else if (io_port_sram_req) begin // @[Reg.scala 28:20]
      stage1_sram_addr_reg <= io_port_sram_addr;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 146:38]
      stage1_sram_phy_addr_reg <= 32'h0; // @[macros.scala 421:45 inst_cache.scala 146:74]
    end else if (stage1_stall_reg) begin
      if (_stage1_sram_phy_addr_reg_T[31:30] == 2'h2) begin
        stage1_sram_phy_addr_reg <= _stage1_sram_phy_addr_reg_T_4;
      end else if (io_tlb_req) begin
        stage1_sram_phy_addr_reg <= io_p_addr_for_tlb;
      end else begin
        stage1_sram_phy_addr_reg <= stage1_sram_addr_reg;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      stage1_sram_cache_reg <= 1'h0; // @[Reg.scala 29:22]
    end else if (io_port_sram_req) begin // @[Reg.scala 28:20]
      stage1_sram_cache_reg <= io_port_sram_cache;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      stage1_sram_req_reg <= 1'h0; // @[Reg.scala 29:22]
    end else if (io_port_sram_req) begin // @[Reg.scala 28:20]
      stage1_sram_req_reg <= io_inst_ready_to_use;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 160:29]
      stage1_sram_valid <= 2'h0;
    end else if (io_port_sram_req) begin // @[inst_cache.scala 153:40]
      stage1_sram_valid <= 2'h3;
    end else if (io_stage1_valid_flush[0]) begin // @[inst_cache.scala 154:12]
      stage1_sram_valid <= 2'h1;
    end else if (io_stage1_valid_flush[1]) begin
      stage1_sram_valid <= 2'h2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 152:27]
      stage1_finished <= 1'h0;
    end else if (io_port_sram_req) begin
      stage1_finished <= 1'h0;
    end else begin
      stage1_finished <= work_state == 4'h7 | work_state == 4'h3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 147:29]
      stage1_exception <= 2'h0;
    end else if (io_port_sram_req) begin
      stage1_exception <= 2'h0;
    end else begin
      stage1_exception <= io_tlb_exception;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 222:29]
      stage2_exception <= 2'h0;
    end else if (stage2_stall) begin // @[inst_cache.scala 222:63]
      stage2_exception <= stage1_exception;
    end else if (io_stage2_flush) begin
      stage2_exception <= 2'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 197:33]
      stage2_sram_addr_reg <= 32'h0;
    end else if (io_stage2_flush) begin // @[inst_cache.scala 197:54]
      stage2_sram_addr_reg <= 32'h0;
    end else if (stage2_stall) begin
      stage2_sram_addr_reg <= stage1_sram_addr_reg;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 206:31]
      stage2_sram_req_reg <= 1'h0;
    end else if (io_stage2_flush) begin // @[inst_cache.scala 206:52]
      stage2_sram_req_reg <= 1'h0;
    end else if (stage2_stall) begin
      stage2_sram_req_reg <= stage1_sram_req_reg;
    end else begin
      stage2_sram_req_reg <= io_port_sram_write_en == 2'h0 & stage2_sram_req_reg;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 210:27]
      stage2_hit0_reg <= 1'h0;
    end else if (io_stage2_flush) begin // @[inst_cache.scala 210:48]
      stage2_hit0_reg <= 1'h0;
    end else if (stage2_stall) begin
      stage2_hit0_reg <= _hit_T_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 229:31]
      stage2_write_en_reg <= 2'h0;
    end else if (io_stage2_flush | io_inst_ready_branch & ~io_inst_buffer_empty) begin // @[inst_cache.scala 229:104]
      stage2_write_en_reg <= 2'h0;
    end else if (stage2_stall) begin
      stage2_write_en_reg <= {{1'd0}, _stage2_write_en_reg_T_17};
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 156:129]
      has_stage2_stall <= 1'h0;
    end else begin
      has_stage2_stall <= (access_work_state == 4'h1 | access_work_state == 4'h4 | stage1_exception != 2'h0) &
        _stage2_stall_T_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 249:28]
      sram_rdata_L_Reg <= 40'h0; // @[inst_cache.scala 238:25 246:{35,84}]
    end else if (has_stage2_stall) begin
      if (_access_work_state_T_8) begin
        sram_rdata_L_Reg <= wait_data_L;
      end else if (_access_work_state_T_23) begin
        if (stage2_hit0_reg) begin
          sram_rdata_L_Reg <= _GEN_522;
        end else begin
          sram_rdata_L_Reg <= _GEN_530;
        end
      end else begin
        sram_rdata_L_Reg <= 40'h0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lru_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  lru_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  lru_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  lru_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  lru_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lru_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  lru_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  lru_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  lru_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  lru_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  lru_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  lru_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  lru_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  lru_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  lru_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  lru_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  lru_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  lru_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  lru_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  lru_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  lru_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  lru_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  lru_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  lru_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  lru_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  lru_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  lru_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  lru_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  lru_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  lru_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  lru_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  lru_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  lru_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  lru_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  lru_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  lru_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  lru_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  lru_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  lru_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  lru_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  lru_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  lru_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  lru_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  lru_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  lru_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  lru_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  lru_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  lru_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  lru_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  lru_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  lru_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  lru_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  lru_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  lru_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  lru_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  lru_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  lru_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  lru_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  lru_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  lru_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  lru_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  lru_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  lru_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  lru_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  lru_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  lru_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  lru_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  lru_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  lru_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  lru_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  lru_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  lru_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  lru_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  lru_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  lru_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  lru_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  lru_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  lru_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  lru_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  lru_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  lru_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  lru_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  lru_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  lru_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  lru_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  lru_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  lru_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  lru_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  lru_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  lru_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  lru_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  lru_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  lru_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  lru_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  lru_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  lru_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  lru_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  lru_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  lru_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  lru_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  lru_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  lru_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  lru_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  lru_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  lru_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  lru_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  lru_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  lru_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  lru_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  lru_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  lru_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  lru_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  lru_112 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  lru_113 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  lru_114 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  lru_115 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  lru_116 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  lru_117 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  lru_118 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  lru_119 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  lru_120 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  lru_121 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  lru_122 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  lru_123 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  lru_124 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  lru_125 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  lru_126 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  lru_127 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  work_state = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  write_counter = _RAND_129[2:0];
  _RAND_130 = {2{`RANDOM}};
  wait_data_L = _RAND_130[39:0];
  _RAND_131 = {1{`RANDOM}};
  stage1_stall_reg = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  stage1_sram_addr_reg = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  stage1_sram_phy_addr_reg = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  stage1_sram_cache_reg = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  stage1_sram_req_reg = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  stage1_sram_valid = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  stage1_finished = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  stage1_exception = _RAND_138[1:0];
  _RAND_139 = {1{`RANDOM}};
  stage2_exception = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  stage2_sram_addr_reg = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  stage2_sram_req_reg = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  stage2_hit0_reg = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  stage2_write_en_reg = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  has_stage2_stall = _RAND_144[0:0];
  _RAND_145 = {2{`RANDOM}};
  sram_rdata_L_Reg = _RAND_145[39:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    lru_0 = 1'h0;
  end
  if (reset) begin
    lru_1 = 1'h0;
  end
  if (reset) begin
    lru_2 = 1'h0;
  end
  if (reset) begin
    lru_3 = 1'h0;
  end
  if (reset) begin
    lru_4 = 1'h0;
  end
  if (reset) begin
    lru_5 = 1'h0;
  end
  if (reset) begin
    lru_6 = 1'h0;
  end
  if (reset) begin
    lru_7 = 1'h0;
  end
  if (reset) begin
    lru_8 = 1'h0;
  end
  if (reset) begin
    lru_9 = 1'h0;
  end
  if (reset) begin
    lru_10 = 1'h0;
  end
  if (reset) begin
    lru_11 = 1'h0;
  end
  if (reset) begin
    lru_12 = 1'h0;
  end
  if (reset) begin
    lru_13 = 1'h0;
  end
  if (reset) begin
    lru_14 = 1'h0;
  end
  if (reset) begin
    lru_15 = 1'h0;
  end
  if (reset) begin
    lru_16 = 1'h0;
  end
  if (reset) begin
    lru_17 = 1'h0;
  end
  if (reset) begin
    lru_18 = 1'h0;
  end
  if (reset) begin
    lru_19 = 1'h0;
  end
  if (reset) begin
    lru_20 = 1'h0;
  end
  if (reset) begin
    lru_21 = 1'h0;
  end
  if (reset) begin
    lru_22 = 1'h0;
  end
  if (reset) begin
    lru_23 = 1'h0;
  end
  if (reset) begin
    lru_24 = 1'h0;
  end
  if (reset) begin
    lru_25 = 1'h0;
  end
  if (reset) begin
    lru_26 = 1'h0;
  end
  if (reset) begin
    lru_27 = 1'h0;
  end
  if (reset) begin
    lru_28 = 1'h0;
  end
  if (reset) begin
    lru_29 = 1'h0;
  end
  if (reset) begin
    lru_30 = 1'h0;
  end
  if (reset) begin
    lru_31 = 1'h0;
  end
  if (reset) begin
    lru_32 = 1'h0;
  end
  if (reset) begin
    lru_33 = 1'h0;
  end
  if (reset) begin
    lru_34 = 1'h0;
  end
  if (reset) begin
    lru_35 = 1'h0;
  end
  if (reset) begin
    lru_36 = 1'h0;
  end
  if (reset) begin
    lru_37 = 1'h0;
  end
  if (reset) begin
    lru_38 = 1'h0;
  end
  if (reset) begin
    lru_39 = 1'h0;
  end
  if (reset) begin
    lru_40 = 1'h0;
  end
  if (reset) begin
    lru_41 = 1'h0;
  end
  if (reset) begin
    lru_42 = 1'h0;
  end
  if (reset) begin
    lru_43 = 1'h0;
  end
  if (reset) begin
    lru_44 = 1'h0;
  end
  if (reset) begin
    lru_45 = 1'h0;
  end
  if (reset) begin
    lru_46 = 1'h0;
  end
  if (reset) begin
    lru_47 = 1'h0;
  end
  if (reset) begin
    lru_48 = 1'h0;
  end
  if (reset) begin
    lru_49 = 1'h0;
  end
  if (reset) begin
    lru_50 = 1'h0;
  end
  if (reset) begin
    lru_51 = 1'h0;
  end
  if (reset) begin
    lru_52 = 1'h0;
  end
  if (reset) begin
    lru_53 = 1'h0;
  end
  if (reset) begin
    lru_54 = 1'h0;
  end
  if (reset) begin
    lru_55 = 1'h0;
  end
  if (reset) begin
    lru_56 = 1'h0;
  end
  if (reset) begin
    lru_57 = 1'h0;
  end
  if (reset) begin
    lru_58 = 1'h0;
  end
  if (reset) begin
    lru_59 = 1'h0;
  end
  if (reset) begin
    lru_60 = 1'h0;
  end
  if (reset) begin
    lru_61 = 1'h0;
  end
  if (reset) begin
    lru_62 = 1'h0;
  end
  if (reset) begin
    lru_63 = 1'h0;
  end
  if (reset) begin
    lru_64 = 1'h0;
  end
  if (reset) begin
    lru_65 = 1'h0;
  end
  if (reset) begin
    lru_66 = 1'h0;
  end
  if (reset) begin
    lru_67 = 1'h0;
  end
  if (reset) begin
    lru_68 = 1'h0;
  end
  if (reset) begin
    lru_69 = 1'h0;
  end
  if (reset) begin
    lru_70 = 1'h0;
  end
  if (reset) begin
    lru_71 = 1'h0;
  end
  if (reset) begin
    lru_72 = 1'h0;
  end
  if (reset) begin
    lru_73 = 1'h0;
  end
  if (reset) begin
    lru_74 = 1'h0;
  end
  if (reset) begin
    lru_75 = 1'h0;
  end
  if (reset) begin
    lru_76 = 1'h0;
  end
  if (reset) begin
    lru_77 = 1'h0;
  end
  if (reset) begin
    lru_78 = 1'h0;
  end
  if (reset) begin
    lru_79 = 1'h0;
  end
  if (reset) begin
    lru_80 = 1'h0;
  end
  if (reset) begin
    lru_81 = 1'h0;
  end
  if (reset) begin
    lru_82 = 1'h0;
  end
  if (reset) begin
    lru_83 = 1'h0;
  end
  if (reset) begin
    lru_84 = 1'h0;
  end
  if (reset) begin
    lru_85 = 1'h0;
  end
  if (reset) begin
    lru_86 = 1'h0;
  end
  if (reset) begin
    lru_87 = 1'h0;
  end
  if (reset) begin
    lru_88 = 1'h0;
  end
  if (reset) begin
    lru_89 = 1'h0;
  end
  if (reset) begin
    lru_90 = 1'h0;
  end
  if (reset) begin
    lru_91 = 1'h0;
  end
  if (reset) begin
    lru_92 = 1'h0;
  end
  if (reset) begin
    lru_93 = 1'h0;
  end
  if (reset) begin
    lru_94 = 1'h0;
  end
  if (reset) begin
    lru_95 = 1'h0;
  end
  if (reset) begin
    lru_96 = 1'h0;
  end
  if (reset) begin
    lru_97 = 1'h0;
  end
  if (reset) begin
    lru_98 = 1'h0;
  end
  if (reset) begin
    lru_99 = 1'h0;
  end
  if (reset) begin
    lru_100 = 1'h0;
  end
  if (reset) begin
    lru_101 = 1'h0;
  end
  if (reset) begin
    lru_102 = 1'h0;
  end
  if (reset) begin
    lru_103 = 1'h0;
  end
  if (reset) begin
    lru_104 = 1'h0;
  end
  if (reset) begin
    lru_105 = 1'h0;
  end
  if (reset) begin
    lru_106 = 1'h0;
  end
  if (reset) begin
    lru_107 = 1'h0;
  end
  if (reset) begin
    lru_108 = 1'h0;
  end
  if (reset) begin
    lru_109 = 1'h0;
  end
  if (reset) begin
    lru_110 = 1'h0;
  end
  if (reset) begin
    lru_111 = 1'h0;
  end
  if (reset) begin
    lru_112 = 1'h0;
  end
  if (reset) begin
    lru_113 = 1'h0;
  end
  if (reset) begin
    lru_114 = 1'h0;
  end
  if (reset) begin
    lru_115 = 1'h0;
  end
  if (reset) begin
    lru_116 = 1'h0;
  end
  if (reset) begin
    lru_117 = 1'h0;
  end
  if (reset) begin
    lru_118 = 1'h0;
  end
  if (reset) begin
    lru_119 = 1'h0;
  end
  if (reset) begin
    lru_120 = 1'h0;
  end
  if (reset) begin
    lru_121 = 1'h0;
  end
  if (reset) begin
    lru_122 = 1'h0;
  end
  if (reset) begin
    lru_123 = 1'h0;
  end
  if (reset) begin
    lru_124 = 1'h0;
  end
  if (reset) begin
    lru_125 = 1'h0;
  end
  if (reset) begin
    lru_126 = 1'h0;
  end
  if (reset) begin
    lru_127 = 1'h0;
  end
  if (reset) begin
    work_state = 4'h1;
  end
  if (reset) begin
    write_counter = 3'h0;
  end
  if (reset) begin
    wait_data_L = 40'h0;
  end
  if (reset) begin
    stage1_stall_reg = 1'h0;
  end
  if (reset) begin
    stage1_sram_addr_reg = 32'h0;
  end
  if (reset) begin
    stage1_sram_phy_addr_reg = 32'h0;
  end
  if (reset) begin
    stage1_sram_cache_reg = 1'h0;
  end
  if (reset) begin
    stage1_sram_req_reg = 1'h0;
  end
  if (reset) begin
    stage1_sram_valid = 2'h0;
  end
  if (reset) begin
    stage1_finished = 1'h0;
  end
  if (reset) begin
    stage1_exception = 2'h0;
  end
  if (reset) begin
    stage2_exception = 2'h0;
  end
  if (reset) begin
    stage2_sram_addr_reg = 32'h0;
  end
  if (reset) begin
    stage2_sram_req_reg = 1'h0;
  end
  if (reset) begin
    stage2_hit0_reg = 1'h0;
  end
  if (reset) begin
    stage2_write_en_reg = 2'h0;
  end
  if (reset) begin
    has_stage2_stall = 1'h0;
  end
  if (reset) begin
    sram_rdata_L_Reg = 40'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module dcache_tag(
  input         clock,
  input         reset,
  input         io_wen,
  input  [20:0] io_wdata,
  input  [31:0] io_raddr,
  input  [31:0] io_waddr,
  output        io_hit,
  output        io_valid,
  output [19:0] io_tag
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
`endif // RANDOMIZE_REG_INIT
  reg [20:0] tag_regs0_0; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_1; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_2; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_3; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_4; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_5; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_6; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_7; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_8; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_9; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_10; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_11; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_12; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_13; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_14; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_15; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_16; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_17; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_18; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_19; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_20; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_21; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_22; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_23; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_24; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_25; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_26; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_27; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_28; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_29; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_30; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_31; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_32; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_33; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_34; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_35; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_36; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_37; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_38; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_39; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_40; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_41; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_42; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_43; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_44; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_45; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_46; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_47; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_48; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_49; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_50; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_51; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_52; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_53; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_54; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_55; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_56; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_57; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_58; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_59; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_60; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_61; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_62; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs0_63; // @[dcache_tag.scala 30:28]
  reg [20:0] tag_regs1_0; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_1; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_2; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_3; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_4; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_5; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_6; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_7; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_8; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_9; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_10; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_11; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_12; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_13; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_14; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_15; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_16; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_17; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_18; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_19; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_20; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_21; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_22; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_23; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_24; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_25; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_26; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_27; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_28; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_29; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_30; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_31; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_32; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_33; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_34; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_35; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_36; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_37; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_38; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_39; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_40; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_41; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_42; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_43; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_44; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_45; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_46; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_47; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_48; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_49; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_50; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_51; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_52; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_53; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_54; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_55; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_56; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_57; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_58; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_59; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_60; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_61; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_62; // @[dcache_tag.scala 31:28]
  reg [20:0] tag_regs1_63; // @[dcache_tag.scala 31:28]
  wire [20:0] _GEN_1 = 6'h1 == io_waddr[11:6] ? tag_regs0_1 : tag_regs0_0; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_2 = 6'h2 == io_waddr[11:6] ? tag_regs0_2 : _GEN_1; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_3 = 6'h3 == io_waddr[11:6] ? tag_regs0_3 : _GEN_2; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_4 = 6'h4 == io_waddr[11:6] ? tag_regs0_4 : _GEN_3; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_5 = 6'h5 == io_waddr[11:6] ? tag_regs0_5 : _GEN_4; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_6 = 6'h6 == io_waddr[11:6] ? tag_regs0_6 : _GEN_5; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_7 = 6'h7 == io_waddr[11:6] ? tag_regs0_7 : _GEN_6; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_8 = 6'h8 == io_waddr[11:6] ? tag_regs0_8 : _GEN_7; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_9 = 6'h9 == io_waddr[11:6] ? tag_regs0_9 : _GEN_8; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_10 = 6'ha == io_waddr[11:6] ? tag_regs0_10 : _GEN_9; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_11 = 6'hb == io_waddr[11:6] ? tag_regs0_11 : _GEN_10; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_12 = 6'hc == io_waddr[11:6] ? tag_regs0_12 : _GEN_11; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_13 = 6'hd == io_waddr[11:6] ? tag_regs0_13 : _GEN_12; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_14 = 6'he == io_waddr[11:6] ? tag_regs0_14 : _GEN_13; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_15 = 6'hf == io_waddr[11:6] ? tag_regs0_15 : _GEN_14; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_16 = 6'h10 == io_waddr[11:6] ? tag_regs0_16 : _GEN_15; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_17 = 6'h11 == io_waddr[11:6] ? tag_regs0_17 : _GEN_16; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_18 = 6'h12 == io_waddr[11:6] ? tag_regs0_18 : _GEN_17; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_19 = 6'h13 == io_waddr[11:6] ? tag_regs0_19 : _GEN_18; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_20 = 6'h14 == io_waddr[11:6] ? tag_regs0_20 : _GEN_19; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_21 = 6'h15 == io_waddr[11:6] ? tag_regs0_21 : _GEN_20; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_22 = 6'h16 == io_waddr[11:6] ? tag_regs0_22 : _GEN_21; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_23 = 6'h17 == io_waddr[11:6] ? tag_regs0_23 : _GEN_22; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_24 = 6'h18 == io_waddr[11:6] ? tag_regs0_24 : _GEN_23; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_25 = 6'h19 == io_waddr[11:6] ? tag_regs0_25 : _GEN_24; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_26 = 6'h1a == io_waddr[11:6] ? tag_regs0_26 : _GEN_25; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_27 = 6'h1b == io_waddr[11:6] ? tag_regs0_27 : _GEN_26; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_28 = 6'h1c == io_waddr[11:6] ? tag_regs0_28 : _GEN_27; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_29 = 6'h1d == io_waddr[11:6] ? tag_regs0_29 : _GEN_28; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_30 = 6'h1e == io_waddr[11:6] ? tag_regs0_30 : _GEN_29; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_31 = 6'h1f == io_waddr[11:6] ? tag_regs0_31 : _GEN_30; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_32 = 6'h20 == io_waddr[11:6] ? tag_regs0_32 : _GEN_31; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_33 = 6'h21 == io_waddr[11:6] ? tag_regs0_33 : _GEN_32; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_34 = 6'h22 == io_waddr[11:6] ? tag_regs0_34 : _GEN_33; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_35 = 6'h23 == io_waddr[11:6] ? tag_regs0_35 : _GEN_34; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_36 = 6'h24 == io_waddr[11:6] ? tag_regs0_36 : _GEN_35; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_37 = 6'h25 == io_waddr[11:6] ? tag_regs0_37 : _GEN_36; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_38 = 6'h26 == io_waddr[11:6] ? tag_regs0_38 : _GEN_37; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_39 = 6'h27 == io_waddr[11:6] ? tag_regs0_39 : _GEN_38; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_40 = 6'h28 == io_waddr[11:6] ? tag_regs0_40 : _GEN_39; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_41 = 6'h29 == io_waddr[11:6] ? tag_regs0_41 : _GEN_40; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_42 = 6'h2a == io_waddr[11:6] ? tag_regs0_42 : _GEN_41; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_43 = 6'h2b == io_waddr[11:6] ? tag_regs0_43 : _GEN_42; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_44 = 6'h2c == io_waddr[11:6] ? tag_regs0_44 : _GEN_43; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_45 = 6'h2d == io_waddr[11:6] ? tag_regs0_45 : _GEN_44; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_46 = 6'h2e == io_waddr[11:6] ? tag_regs0_46 : _GEN_45; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_47 = 6'h2f == io_waddr[11:6] ? tag_regs0_47 : _GEN_46; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_48 = 6'h30 == io_waddr[11:6] ? tag_regs0_48 : _GEN_47; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_49 = 6'h31 == io_waddr[11:6] ? tag_regs0_49 : _GEN_48; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_50 = 6'h32 == io_waddr[11:6] ? tag_regs0_50 : _GEN_49; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_51 = 6'h33 == io_waddr[11:6] ? tag_regs0_51 : _GEN_50; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_52 = 6'h34 == io_waddr[11:6] ? tag_regs0_52 : _GEN_51; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_53 = 6'h35 == io_waddr[11:6] ? tag_regs0_53 : _GEN_52; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_54 = 6'h36 == io_waddr[11:6] ? tag_regs0_54 : _GEN_53; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_55 = 6'h37 == io_waddr[11:6] ? tag_regs0_55 : _GEN_54; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_56 = 6'h38 == io_waddr[11:6] ? tag_regs0_56 : _GEN_55; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_57 = 6'h39 == io_waddr[11:6] ? tag_regs0_57 : _GEN_56; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_58 = 6'h3a == io_waddr[11:6] ? tag_regs0_58 : _GEN_57; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_59 = 6'h3b == io_waddr[11:6] ? tag_regs0_59 : _GEN_58; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_60 = 6'h3c == io_waddr[11:6] ? tag_regs0_60 : _GEN_59; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_61 = 6'h3d == io_waddr[11:6] ? tag_regs0_61 : _GEN_60; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_62 = 6'h3e == io_waddr[11:6] ? tag_regs0_62 : _GEN_61; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_63 = 6'h3f == io_waddr[11:6] ? tag_regs0_63 : _GEN_62; // @[dcache_tag.scala 34:{37,37}]
  wire [20:0] _GEN_129 = 6'h1 == io_waddr[11:6] ? tag_regs1_1 : tag_regs1_0; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_130 = 6'h2 == io_waddr[11:6] ? tag_regs1_2 : _GEN_129; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_131 = 6'h3 == io_waddr[11:6] ? tag_regs1_3 : _GEN_130; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_132 = 6'h4 == io_waddr[11:6] ? tag_regs1_4 : _GEN_131; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_133 = 6'h5 == io_waddr[11:6] ? tag_regs1_5 : _GEN_132; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_134 = 6'h6 == io_waddr[11:6] ? tag_regs1_6 : _GEN_133; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_135 = 6'h7 == io_waddr[11:6] ? tag_regs1_7 : _GEN_134; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_136 = 6'h8 == io_waddr[11:6] ? tag_regs1_8 : _GEN_135; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_137 = 6'h9 == io_waddr[11:6] ? tag_regs1_9 : _GEN_136; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_138 = 6'ha == io_waddr[11:6] ? tag_regs1_10 : _GEN_137; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_139 = 6'hb == io_waddr[11:6] ? tag_regs1_11 : _GEN_138; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_140 = 6'hc == io_waddr[11:6] ? tag_regs1_12 : _GEN_139; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_141 = 6'hd == io_waddr[11:6] ? tag_regs1_13 : _GEN_140; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_142 = 6'he == io_waddr[11:6] ? tag_regs1_14 : _GEN_141; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_143 = 6'hf == io_waddr[11:6] ? tag_regs1_15 : _GEN_142; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_144 = 6'h10 == io_waddr[11:6] ? tag_regs1_16 : _GEN_143; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_145 = 6'h11 == io_waddr[11:6] ? tag_regs1_17 : _GEN_144; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_146 = 6'h12 == io_waddr[11:6] ? tag_regs1_18 : _GEN_145; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_147 = 6'h13 == io_waddr[11:6] ? tag_regs1_19 : _GEN_146; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_148 = 6'h14 == io_waddr[11:6] ? tag_regs1_20 : _GEN_147; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_149 = 6'h15 == io_waddr[11:6] ? tag_regs1_21 : _GEN_148; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_150 = 6'h16 == io_waddr[11:6] ? tag_regs1_22 : _GEN_149; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_151 = 6'h17 == io_waddr[11:6] ? tag_regs1_23 : _GEN_150; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_152 = 6'h18 == io_waddr[11:6] ? tag_regs1_24 : _GEN_151; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_153 = 6'h19 == io_waddr[11:6] ? tag_regs1_25 : _GEN_152; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_154 = 6'h1a == io_waddr[11:6] ? tag_regs1_26 : _GEN_153; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_155 = 6'h1b == io_waddr[11:6] ? tag_regs1_27 : _GEN_154; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_156 = 6'h1c == io_waddr[11:6] ? tag_regs1_28 : _GEN_155; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_157 = 6'h1d == io_waddr[11:6] ? tag_regs1_29 : _GEN_156; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_158 = 6'h1e == io_waddr[11:6] ? tag_regs1_30 : _GEN_157; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_159 = 6'h1f == io_waddr[11:6] ? tag_regs1_31 : _GEN_158; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_160 = 6'h20 == io_waddr[11:6] ? tag_regs1_32 : _GEN_159; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_161 = 6'h21 == io_waddr[11:6] ? tag_regs1_33 : _GEN_160; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_162 = 6'h22 == io_waddr[11:6] ? tag_regs1_34 : _GEN_161; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_163 = 6'h23 == io_waddr[11:6] ? tag_regs1_35 : _GEN_162; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_164 = 6'h24 == io_waddr[11:6] ? tag_regs1_36 : _GEN_163; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_165 = 6'h25 == io_waddr[11:6] ? tag_regs1_37 : _GEN_164; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_166 = 6'h26 == io_waddr[11:6] ? tag_regs1_38 : _GEN_165; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_167 = 6'h27 == io_waddr[11:6] ? tag_regs1_39 : _GEN_166; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_168 = 6'h28 == io_waddr[11:6] ? tag_regs1_40 : _GEN_167; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_169 = 6'h29 == io_waddr[11:6] ? tag_regs1_41 : _GEN_168; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_170 = 6'h2a == io_waddr[11:6] ? tag_regs1_42 : _GEN_169; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_171 = 6'h2b == io_waddr[11:6] ? tag_regs1_43 : _GEN_170; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_172 = 6'h2c == io_waddr[11:6] ? tag_regs1_44 : _GEN_171; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_173 = 6'h2d == io_waddr[11:6] ? tag_regs1_45 : _GEN_172; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_174 = 6'h2e == io_waddr[11:6] ? tag_regs1_46 : _GEN_173; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_175 = 6'h2f == io_waddr[11:6] ? tag_regs1_47 : _GEN_174; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_176 = 6'h30 == io_waddr[11:6] ? tag_regs1_48 : _GEN_175; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_177 = 6'h31 == io_waddr[11:6] ? tag_regs1_49 : _GEN_176; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_178 = 6'h32 == io_waddr[11:6] ? tag_regs1_50 : _GEN_177; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_179 = 6'h33 == io_waddr[11:6] ? tag_regs1_51 : _GEN_178; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_180 = 6'h34 == io_waddr[11:6] ? tag_regs1_52 : _GEN_179; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_181 = 6'h35 == io_waddr[11:6] ? tag_regs1_53 : _GEN_180; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_182 = 6'h36 == io_waddr[11:6] ? tag_regs1_54 : _GEN_181; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_183 = 6'h37 == io_waddr[11:6] ? tag_regs1_55 : _GEN_182; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_184 = 6'h38 == io_waddr[11:6] ? tag_regs1_56 : _GEN_183; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_185 = 6'h39 == io_waddr[11:6] ? tag_regs1_57 : _GEN_184; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_186 = 6'h3a == io_waddr[11:6] ? tag_regs1_58 : _GEN_185; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_187 = 6'h3b == io_waddr[11:6] ? tag_regs1_59 : _GEN_186; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_188 = 6'h3c == io_waddr[11:6] ? tag_regs1_60 : _GEN_187; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_189 = 6'h3d == io_waddr[11:6] ? tag_regs1_61 : _GEN_188; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_190 = 6'h3e == io_waddr[11:6] ? tag_regs1_62 : _GEN_189; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_191 = 6'h3f == io_waddr[11:6] ? tag_regs1_63 : _GEN_190; // @[dcache_tag.scala 35:{37,37}]
  wire [20:0] _GEN_385 = 6'h1 == io_raddr[11:6] ? tag_regs1_1 : tag_regs1_0; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_386 = 6'h2 == io_raddr[11:6] ? tag_regs1_2 : _GEN_385; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_387 = 6'h3 == io_raddr[11:6] ? tag_regs1_3 : _GEN_386; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_388 = 6'h4 == io_raddr[11:6] ? tag_regs1_4 : _GEN_387; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_389 = 6'h5 == io_raddr[11:6] ? tag_regs1_5 : _GEN_388; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_390 = 6'h6 == io_raddr[11:6] ? tag_regs1_6 : _GEN_389; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_391 = 6'h7 == io_raddr[11:6] ? tag_regs1_7 : _GEN_390; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_392 = 6'h8 == io_raddr[11:6] ? tag_regs1_8 : _GEN_391; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_393 = 6'h9 == io_raddr[11:6] ? tag_regs1_9 : _GEN_392; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_394 = 6'ha == io_raddr[11:6] ? tag_regs1_10 : _GEN_393; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_395 = 6'hb == io_raddr[11:6] ? tag_regs1_11 : _GEN_394; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_396 = 6'hc == io_raddr[11:6] ? tag_regs1_12 : _GEN_395; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_397 = 6'hd == io_raddr[11:6] ? tag_regs1_13 : _GEN_396; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_398 = 6'he == io_raddr[11:6] ? tag_regs1_14 : _GEN_397; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_399 = 6'hf == io_raddr[11:6] ? tag_regs1_15 : _GEN_398; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_400 = 6'h10 == io_raddr[11:6] ? tag_regs1_16 : _GEN_399; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_401 = 6'h11 == io_raddr[11:6] ? tag_regs1_17 : _GEN_400; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_402 = 6'h12 == io_raddr[11:6] ? tag_regs1_18 : _GEN_401; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_403 = 6'h13 == io_raddr[11:6] ? tag_regs1_19 : _GEN_402; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_404 = 6'h14 == io_raddr[11:6] ? tag_regs1_20 : _GEN_403; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_405 = 6'h15 == io_raddr[11:6] ? tag_regs1_21 : _GEN_404; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_406 = 6'h16 == io_raddr[11:6] ? tag_regs1_22 : _GEN_405; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_407 = 6'h17 == io_raddr[11:6] ? tag_regs1_23 : _GEN_406; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_408 = 6'h18 == io_raddr[11:6] ? tag_regs1_24 : _GEN_407; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_409 = 6'h19 == io_raddr[11:6] ? tag_regs1_25 : _GEN_408; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_410 = 6'h1a == io_raddr[11:6] ? tag_regs1_26 : _GEN_409; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_411 = 6'h1b == io_raddr[11:6] ? tag_regs1_27 : _GEN_410; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_412 = 6'h1c == io_raddr[11:6] ? tag_regs1_28 : _GEN_411; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_413 = 6'h1d == io_raddr[11:6] ? tag_regs1_29 : _GEN_412; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_414 = 6'h1e == io_raddr[11:6] ? tag_regs1_30 : _GEN_413; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_415 = 6'h1f == io_raddr[11:6] ? tag_regs1_31 : _GEN_414; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_416 = 6'h20 == io_raddr[11:6] ? tag_regs1_32 : _GEN_415; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_417 = 6'h21 == io_raddr[11:6] ? tag_regs1_33 : _GEN_416; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_418 = 6'h22 == io_raddr[11:6] ? tag_regs1_34 : _GEN_417; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_419 = 6'h23 == io_raddr[11:6] ? tag_regs1_35 : _GEN_418; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_420 = 6'h24 == io_raddr[11:6] ? tag_regs1_36 : _GEN_419; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_421 = 6'h25 == io_raddr[11:6] ? tag_regs1_37 : _GEN_420; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_422 = 6'h26 == io_raddr[11:6] ? tag_regs1_38 : _GEN_421; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_423 = 6'h27 == io_raddr[11:6] ? tag_regs1_39 : _GEN_422; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_424 = 6'h28 == io_raddr[11:6] ? tag_regs1_40 : _GEN_423; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_425 = 6'h29 == io_raddr[11:6] ? tag_regs1_41 : _GEN_424; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_426 = 6'h2a == io_raddr[11:6] ? tag_regs1_42 : _GEN_425; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_427 = 6'h2b == io_raddr[11:6] ? tag_regs1_43 : _GEN_426; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_428 = 6'h2c == io_raddr[11:6] ? tag_regs1_44 : _GEN_427; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_429 = 6'h2d == io_raddr[11:6] ? tag_regs1_45 : _GEN_428; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_430 = 6'h2e == io_raddr[11:6] ? tag_regs1_46 : _GEN_429; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_431 = 6'h2f == io_raddr[11:6] ? tag_regs1_47 : _GEN_430; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_432 = 6'h30 == io_raddr[11:6] ? tag_regs1_48 : _GEN_431; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_433 = 6'h31 == io_raddr[11:6] ? tag_regs1_49 : _GEN_432; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_434 = 6'h32 == io_raddr[11:6] ? tag_regs1_50 : _GEN_433; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_435 = 6'h33 == io_raddr[11:6] ? tag_regs1_51 : _GEN_434; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_436 = 6'h34 == io_raddr[11:6] ? tag_regs1_52 : _GEN_435; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_437 = 6'h35 == io_raddr[11:6] ? tag_regs1_53 : _GEN_436; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_438 = 6'h36 == io_raddr[11:6] ? tag_regs1_54 : _GEN_437; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_439 = 6'h37 == io_raddr[11:6] ? tag_regs1_55 : _GEN_438; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_440 = 6'h38 == io_raddr[11:6] ? tag_regs1_56 : _GEN_439; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_441 = 6'h39 == io_raddr[11:6] ? tag_regs1_57 : _GEN_440; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_442 = 6'h3a == io_raddr[11:6] ? tag_regs1_58 : _GEN_441; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_443 = 6'h3b == io_raddr[11:6] ? tag_regs1_59 : _GEN_442; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_444 = 6'h3c == io_raddr[11:6] ? tag_regs1_60 : _GEN_443; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_445 = 6'h3d == io_raddr[11:6] ? tag_regs1_61 : _GEN_444; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_446 = 6'h3e == io_raddr[11:6] ? tag_regs1_62 : _GEN_445; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_447 = 6'h3f == io_raddr[11:6] ? tag_regs1_63 : _GEN_446; // @[dcache_tag.scala 44:{44,44}]
  wire [20:0] _GEN_449 = 6'h1 == io_raddr[11:6] ? tag_regs0_1 : tag_regs0_0; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_450 = 6'h2 == io_raddr[11:6] ? tag_regs0_2 : _GEN_449; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_451 = 6'h3 == io_raddr[11:6] ? tag_regs0_3 : _GEN_450; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_452 = 6'h4 == io_raddr[11:6] ? tag_regs0_4 : _GEN_451; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_453 = 6'h5 == io_raddr[11:6] ? tag_regs0_5 : _GEN_452; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_454 = 6'h6 == io_raddr[11:6] ? tag_regs0_6 : _GEN_453; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_455 = 6'h7 == io_raddr[11:6] ? tag_regs0_7 : _GEN_454; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_456 = 6'h8 == io_raddr[11:6] ? tag_regs0_8 : _GEN_455; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_457 = 6'h9 == io_raddr[11:6] ? tag_regs0_9 : _GEN_456; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_458 = 6'ha == io_raddr[11:6] ? tag_regs0_10 : _GEN_457; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_459 = 6'hb == io_raddr[11:6] ? tag_regs0_11 : _GEN_458; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_460 = 6'hc == io_raddr[11:6] ? tag_regs0_12 : _GEN_459; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_461 = 6'hd == io_raddr[11:6] ? tag_regs0_13 : _GEN_460; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_462 = 6'he == io_raddr[11:6] ? tag_regs0_14 : _GEN_461; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_463 = 6'hf == io_raddr[11:6] ? tag_regs0_15 : _GEN_462; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_464 = 6'h10 == io_raddr[11:6] ? tag_regs0_16 : _GEN_463; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_465 = 6'h11 == io_raddr[11:6] ? tag_regs0_17 : _GEN_464; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_466 = 6'h12 == io_raddr[11:6] ? tag_regs0_18 : _GEN_465; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_467 = 6'h13 == io_raddr[11:6] ? tag_regs0_19 : _GEN_466; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_468 = 6'h14 == io_raddr[11:6] ? tag_regs0_20 : _GEN_467; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_469 = 6'h15 == io_raddr[11:6] ? tag_regs0_21 : _GEN_468; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_470 = 6'h16 == io_raddr[11:6] ? tag_regs0_22 : _GEN_469; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_471 = 6'h17 == io_raddr[11:6] ? tag_regs0_23 : _GEN_470; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_472 = 6'h18 == io_raddr[11:6] ? tag_regs0_24 : _GEN_471; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_473 = 6'h19 == io_raddr[11:6] ? tag_regs0_25 : _GEN_472; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_474 = 6'h1a == io_raddr[11:6] ? tag_regs0_26 : _GEN_473; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_475 = 6'h1b == io_raddr[11:6] ? tag_regs0_27 : _GEN_474; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_476 = 6'h1c == io_raddr[11:6] ? tag_regs0_28 : _GEN_475; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_477 = 6'h1d == io_raddr[11:6] ? tag_regs0_29 : _GEN_476; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_478 = 6'h1e == io_raddr[11:6] ? tag_regs0_30 : _GEN_477; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_479 = 6'h1f == io_raddr[11:6] ? tag_regs0_31 : _GEN_478; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_480 = 6'h20 == io_raddr[11:6] ? tag_regs0_32 : _GEN_479; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_481 = 6'h21 == io_raddr[11:6] ? tag_regs0_33 : _GEN_480; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_482 = 6'h22 == io_raddr[11:6] ? tag_regs0_34 : _GEN_481; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_483 = 6'h23 == io_raddr[11:6] ? tag_regs0_35 : _GEN_482; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_484 = 6'h24 == io_raddr[11:6] ? tag_regs0_36 : _GEN_483; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_485 = 6'h25 == io_raddr[11:6] ? tag_regs0_37 : _GEN_484; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_486 = 6'h26 == io_raddr[11:6] ? tag_regs0_38 : _GEN_485; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_487 = 6'h27 == io_raddr[11:6] ? tag_regs0_39 : _GEN_486; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_488 = 6'h28 == io_raddr[11:6] ? tag_regs0_40 : _GEN_487; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_489 = 6'h29 == io_raddr[11:6] ? tag_regs0_41 : _GEN_488; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_490 = 6'h2a == io_raddr[11:6] ? tag_regs0_42 : _GEN_489; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_491 = 6'h2b == io_raddr[11:6] ? tag_regs0_43 : _GEN_490; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_492 = 6'h2c == io_raddr[11:6] ? tag_regs0_44 : _GEN_491; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_493 = 6'h2d == io_raddr[11:6] ? tag_regs0_45 : _GEN_492; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_494 = 6'h2e == io_raddr[11:6] ? tag_regs0_46 : _GEN_493; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_495 = 6'h2f == io_raddr[11:6] ? tag_regs0_47 : _GEN_494; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_496 = 6'h30 == io_raddr[11:6] ? tag_regs0_48 : _GEN_495; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_497 = 6'h31 == io_raddr[11:6] ? tag_regs0_49 : _GEN_496; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_498 = 6'h32 == io_raddr[11:6] ? tag_regs0_50 : _GEN_497; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_499 = 6'h33 == io_raddr[11:6] ? tag_regs0_51 : _GEN_498; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_500 = 6'h34 == io_raddr[11:6] ? tag_regs0_52 : _GEN_499; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_501 = 6'h35 == io_raddr[11:6] ? tag_regs0_53 : _GEN_500; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_502 = 6'h36 == io_raddr[11:6] ? tag_regs0_54 : _GEN_501; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_503 = 6'h37 == io_raddr[11:6] ? tag_regs0_55 : _GEN_502; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_504 = 6'h38 == io_raddr[11:6] ? tag_regs0_56 : _GEN_503; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_505 = 6'h39 == io_raddr[11:6] ? tag_regs0_57 : _GEN_504; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_506 = 6'h3a == io_raddr[11:6] ? tag_regs0_58 : _GEN_505; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_507 = 6'h3b == io_raddr[11:6] ? tag_regs0_59 : _GEN_506; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_508 = 6'h3c == io_raddr[11:6] ? tag_regs0_60 : _GEN_507; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_509 = 6'h3d == io_raddr[11:6] ? tag_regs0_61 : _GEN_508; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_510 = 6'h3e == io_raddr[11:6] ? tag_regs0_62 : _GEN_509; // @[dcache_tag.scala 44:{60,60}]
  wire [20:0] _GEN_511 = 6'h3f == io_raddr[11:6] ? tag_regs0_63 : _GEN_510; // @[dcache_tag.scala 44:{60,60}]
  assign io_hit = io_raddr[5] & _GEN_447[19:0] == io_raddr[31:12] | ~io_raddr[5] & _GEN_511[19:0] == io_raddr[31:12]; // @[dcache_tag.scala 45:70]
  assign io_valid = io_raddr[5] ? _GEN_447[20] : _GEN_511[20]; // @[dcache_tag.scala 44:20]
  assign io_tag = io_waddr[5] ? _GEN_191[19:0] : _GEN_63[19:0]; // @[dcache_tag.scala 42:18]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_0 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h0 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_0 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_0 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_0 <= tag_regs0_62;
      end else begin
        tag_regs0_0 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_1 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h1 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_1 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_1 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_1 <= tag_regs0_62;
      end else begin
        tag_regs0_1 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_2 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h2 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_2 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_2 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_2 <= tag_regs0_62;
      end else begin
        tag_regs0_2 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_3 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h3 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_3 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_3 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_3 <= tag_regs0_62;
      end else begin
        tag_regs0_3 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_4 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h4 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_4 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_4 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_4 <= tag_regs0_62;
      end else begin
        tag_regs0_4 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_5 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h5 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_5 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_5 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_5 <= tag_regs0_62;
      end else begin
        tag_regs0_5 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_6 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h6 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_6 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_6 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_6 <= tag_regs0_62;
      end else begin
        tag_regs0_6 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_7 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h7 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_7 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_7 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_7 <= tag_regs0_62;
      end else begin
        tag_regs0_7 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_8 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h8 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_8 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_8 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_8 <= tag_regs0_62;
      end else begin
        tag_regs0_8 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_9 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h9 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_9 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_9 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_9 <= tag_regs0_62;
      end else begin
        tag_regs0_9 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_10 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'ha == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_10 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_10 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_10 <= tag_regs0_62;
      end else begin
        tag_regs0_10 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_11 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'hb == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_11 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_11 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_11 <= tag_regs0_62;
      end else begin
        tag_regs0_11 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_12 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'hc == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_12 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_12 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_12 <= tag_regs0_62;
      end else begin
        tag_regs0_12 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_13 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'hd == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_13 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_13 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_13 <= tag_regs0_62;
      end else begin
        tag_regs0_13 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_14 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'he == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_14 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_14 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_14 <= tag_regs0_62;
      end else begin
        tag_regs0_14 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_15 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'hf == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_15 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_15 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_15 <= tag_regs0_62;
      end else begin
        tag_regs0_15 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_16 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h10 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_16 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_16 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_16 <= tag_regs0_62;
      end else begin
        tag_regs0_16 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_17 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h11 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_17 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_17 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_17 <= tag_regs0_62;
      end else begin
        tag_regs0_17 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_18 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h12 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_18 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_18 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_18 <= tag_regs0_62;
      end else begin
        tag_regs0_18 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_19 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h13 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_19 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_19 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_19 <= tag_regs0_62;
      end else begin
        tag_regs0_19 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_20 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h14 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_20 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_20 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_20 <= tag_regs0_62;
      end else begin
        tag_regs0_20 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_21 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h15 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_21 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_21 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_21 <= tag_regs0_62;
      end else begin
        tag_regs0_21 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_22 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h16 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_22 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_22 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_22 <= tag_regs0_62;
      end else begin
        tag_regs0_22 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_23 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h17 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_23 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_23 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_23 <= tag_regs0_62;
      end else begin
        tag_regs0_23 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_24 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h18 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_24 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_24 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_24 <= tag_regs0_62;
      end else begin
        tag_regs0_24 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_25 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h19 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_25 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_25 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_25 <= tag_regs0_62;
      end else begin
        tag_regs0_25 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_26 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h1a == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_26 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_26 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_26 <= tag_regs0_62;
      end else begin
        tag_regs0_26 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_27 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h1b == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_27 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_27 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_27 <= tag_regs0_62;
      end else begin
        tag_regs0_27 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_28 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h1c == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_28 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_28 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_28 <= tag_regs0_62;
      end else begin
        tag_regs0_28 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_29 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h1d == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_29 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_29 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_29 <= tag_regs0_62;
      end else begin
        tag_regs0_29 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_30 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h1e == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_30 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_30 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_30 <= tag_regs0_62;
      end else begin
        tag_regs0_30 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_31 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h1f == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_31 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_31 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_31 <= tag_regs0_62;
      end else begin
        tag_regs0_31 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_32 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h20 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_32 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_32 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_32 <= tag_regs0_62;
      end else begin
        tag_regs0_32 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_33 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h21 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_33 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_33 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_33 <= tag_regs0_62;
      end else begin
        tag_regs0_33 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_34 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h22 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_34 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_34 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_34 <= tag_regs0_62;
      end else begin
        tag_regs0_34 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_35 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h23 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_35 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_35 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_35 <= tag_regs0_62;
      end else begin
        tag_regs0_35 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_36 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h24 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_36 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_36 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_36 <= tag_regs0_62;
      end else begin
        tag_regs0_36 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_37 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h25 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_37 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_37 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_37 <= tag_regs0_62;
      end else begin
        tag_regs0_37 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_38 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h26 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_38 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_38 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_38 <= tag_regs0_62;
      end else begin
        tag_regs0_38 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_39 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h27 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_39 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_39 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_39 <= tag_regs0_62;
      end else begin
        tag_regs0_39 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_40 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h28 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_40 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_40 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_40 <= tag_regs0_62;
      end else begin
        tag_regs0_40 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_41 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h29 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_41 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_41 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_41 <= tag_regs0_62;
      end else begin
        tag_regs0_41 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_42 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h2a == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_42 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_42 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_42 <= tag_regs0_62;
      end else begin
        tag_regs0_42 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_43 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h2b == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_43 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_43 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_43 <= tag_regs0_62;
      end else begin
        tag_regs0_43 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_44 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h2c == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_44 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_44 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_44 <= tag_regs0_62;
      end else begin
        tag_regs0_44 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_45 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h2d == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_45 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_45 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_45 <= tag_regs0_62;
      end else begin
        tag_regs0_45 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_46 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h2e == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_46 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_46 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_46 <= tag_regs0_62;
      end else begin
        tag_regs0_46 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_47 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h2f == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_47 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_47 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_47 <= tag_regs0_62;
      end else begin
        tag_regs0_47 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_48 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h30 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_48 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_48 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_48 <= tag_regs0_62;
      end else begin
        tag_regs0_48 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_49 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h31 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_49 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_49 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_49 <= tag_regs0_62;
      end else begin
        tag_regs0_49 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_50 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h32 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_50 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_50 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_50 <= tag_regs0_62;
      end else begin
        tag_regs0_50 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_51 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h33 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_51 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_51 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_51 <= tag_regs0_62;
      end else begin
        tag_regs0_51 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_52 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h34 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_52 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_52 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_52 <= tag_regs0_62;
      end else begin
        tag_regs0_52 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_53 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h35 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_53 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_53 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_53 <= tag_regs0_62;
      end else begin
        tag_regs0_53 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_54 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h36 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_54 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_54 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_54 <= tag_regs0_62;
      end else begin
        tag_regs0_54 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_55 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h37 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_55 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_55 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_55 <= tag_regs0_62;
      end else begin
        tag_regs0_55 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_56 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h38 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_56 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_56 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_56 <= tag_regs0_62;
      end else begin
        tag_regs0_56 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_57 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h39 == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_57 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_57 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_57 <= tag_regs0_62;
      end else begin
        tag_regs0_57 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_58 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h3a == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_58 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_58 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_58 <= tag_regs0_62;
      end else begin
        tag_regs0_58 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_59 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h3b == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_59 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_59 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_59 <= tag_regs0_62;
      end else begin
        tag_regs0_59 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_60 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h3c == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_60 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_60 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_60 <= tag_regs0_62;
      end else begin
        tag_regs0_60 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_61 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h3d == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_61 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_61 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs0_61 <= tag_regs0_62;
      end else begin
        tag_regs0_61 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_62 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h3e == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_62 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs0_62 <= tag_regs0_63;
      end else if (!(6'h3e == io_waddr[11:6])) begin
        tag_regs0_62 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 34:31]
      tag_regs0_63 <= 21'h0; // @[dcache_tag.scala 34:{37,37,37,37,37}]
    end else if (6'h3f == io_waddr[11:6]) begin // @[dcache_tag.scala 30:28]
      if (io_wen & ~io_waddr[5]) begin
        tag_regs0_63 <= io_wdata;
      end else if (!(6'h3f == io_waddr[11:6])) begin
        if (6'h3e == io_waddr[11:6]) begin
          tag_regs0_63 <= tag_regs0_62;
        end else begin
          tag_regs0_63 <= _GEN_61;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_0 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h0 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_0 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_0 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_0 <= tag_regs1_62;
      end else begin
        tag_regs1_0 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_1 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h1 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_1 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_1 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_1 <= tag_regs1_62;
      end else begin
        tag_regs1_1 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_2 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h2 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_2 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_2 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_2 <= tag_regs1_62;
      end else begin
        tag_regs1_2 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_3 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h3 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_3 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_3 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_3 <= tag_regs1_62;
      end else begin
        tag_regs1_3 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_4 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h4 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_4 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_4 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_4 <= tag_regs1_62;
      end else begin
        tag_regs1_4 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_5 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h5 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_5 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_5 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_5 <= tag_regs1_62;
      end else begin
        tag_regs1_5 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_6 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h6 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_6 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_6 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_6 <= tag_regs1_62;
      end else begin
        tag_regs1_6 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_7 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h7 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_7 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_7 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_7 <= tag_regs1_62;
      end else begin
        tag_regs1_7 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_8 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h8 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_8 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_8 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_8 <= tag_regs1_62;
      end else begin
        tag_regs1_8 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_9 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h9 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_9 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_9 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_9 <= tag_regs1_62;
      end else begin
        tag_regs1_9 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_10 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'ha == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_10 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_10 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_10 <= tag_regs1_62;
      end else begin
        tag_regs1_10 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_11 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'hb == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_11 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_11 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_11 <= tag_regs1_62;
      end else begin
        tag_regs1_11 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_12 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'hc == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_12 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_12 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_12 <= tag_regs1_62;
      end else begin
        tag_regs1_12 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_13 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'hd == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_13 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_13 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_13 <= tag_regs1_62;
      end else begin
        tag_regs1_13 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_14 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'he == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_14 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_14 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_14 <= tag_regs1_62;
      end else begin
        tag_regs1_14 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_15 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'hf == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_15 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_15 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_15 <= tag_regs1_62;
      end else begin
        tag_regs1_15 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_16 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h10 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_16 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_16 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_16 <= tag_regs1_62;
      end else begin
        tag_regs1_16 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_17 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h11 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_17 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_17 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_17 <= tag_regs1_62;
      end else begin
        tag_regs1_17 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_18 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h12 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_18 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_18 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_18 <= tag_regs1_62;
      end else begin
        tag_regs1_18 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_19 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h13 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_19 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_19 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_19 <= tag_regs1_62;
      end else begin
        tag_regs1_19 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_20 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h14 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_20 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_20 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_20 <= tag_regs1_62;
      end else begin
        tag_regs1_20 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_21 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h15 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_21 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_21 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_21 <= tag_regs1_62;
      end else begin
        tag_regs1_21 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_22 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h16 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_22 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_22 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_22 <= tag_regs1_62;
      end else begin
        tag_regs1_22 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_23 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h17 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_23 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_23 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_23 <= tag_regs1_62;
      end else begin
        tag_regs1_23 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_24 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h18 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_24 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_24 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_24 <= tag_regs1_62;
      end else begin
        tag_regs1_24 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_25 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h19 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_25 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_25 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_25 <= tag_regs1_62;
      end else begin
        tag_regs1_25 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_26 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h1a == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_26 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_26 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_26 <= tag_regs1_62;
      end else begin
        tag_regs1_26 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_27 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h1b == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_27 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_27 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_27 <= tag_regs1_62;
      end else begin
        tag_regs1_27 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_28 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h1c == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_28 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_28 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_28 <= tag_regs1_62;
      end else begin
        tag_regs1_28 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_29 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h1d == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_29 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_29 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_29 <= tag_regs1_62;
      end else begin
        tag_regs1_29 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_30 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h1e == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_30 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_30 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_30 <= tag_regs1_62;
      end else begin
        tag_regs1_30 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_31 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h1f == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_31 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_31 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_31 <= tag_regs1_62;
      end else begin
        tag_regs1_31 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_32 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h20 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_32 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_32 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_32 <= tag_regs1_62;
      end else begin
        tag_regs1_32 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_33 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h21 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_33 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_33 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_33 <= tag_regs1_62;
      end else begin
        tag_regs1_33 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_34 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h22 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_34 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_34 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_34 <= tag_regs1_62;
      end else begin
        tag_regs1_34 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_35 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h23 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_35 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_35 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_35 <= tag_regs1_62;
      end else begin
        tag_regs1_35 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_36 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h24 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_36 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_36 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_36 <= tag_regs1_62;
      end else begin
        tag_regs1_36 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_37 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h25 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_37 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_37 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_37 <= tag_regs1_62;
      end else begin
        tag_regs1_37 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_38 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h26 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_38 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_38 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_38 <= tag_regs1_62;
      end else begin
        tag_regs1_38 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_39 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h27 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_39 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_39 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_39 <= tag_regs1_62;
      end else begin
        tag_regs1_39 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_40 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h28 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_40 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_40 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_40 <= tag_regs1_62;
      end else begin
        tag_regs1_40 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_41 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h29 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_41 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_41 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_41 <= tag_regs1_62;
      end else begin
        tag_regs1_41 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_42 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h2a == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_42 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_42 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_42 <= tag_regs1_62;
      end else begin
        tag_regs1_42 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_43 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h2b == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_43 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_43 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_43 <= tag_regs1_62;
      end else begin
        tag_regs1_43 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_44 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h2c == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_44 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_44 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_44 <= tag_regs1_62;
      end else begin
        tag_regs1_44 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_45 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h2d == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_45 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_45 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_45 <= tag_regs1_62;
      end else begin
        tag_regs1_45 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_46 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h2e == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_46 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_46 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_46 <= tag_regs1_62;
      end else begin
        tag_regs1_46 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_47 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h2f == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_47 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_47 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_47 <= tag_regs1_62;
      end else begin
        tag_regs1_47 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_48 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h30 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_48 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_48 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_48 <= tag_regs1_62;
      end else begin
        tag_regs1_48 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_49 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h31 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_49 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_49 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_49 <= tag_regs1_62;
      end else begin
        tag_regs1_49 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_50 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h32 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_50 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_50 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_50 <= tag_regs1_62;
      end else begin
        tag_regs1_50 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_51 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h33 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_51 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_51 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_51 <= tag_regs1_62;
      end else begin
        tag_regs1_51 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_52 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h34 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_52 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_52 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_52 <= tag_regs1_62;
      end else begin
        tag_regs1_52 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_53 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h35 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_53 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_53 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_53 <= tag_regs1_62;
      end else begin
        tag_regs1_53 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_54 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h36 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_54 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_54 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_54 <= tag_regs1_62;
      end else begin
        tag_regs1_54 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_55 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h37 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_55 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_55 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_55 <= tag_regs1_62;
      end else begin
        tag_regs1_55 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_56 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h38 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_56 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_56 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_56 <= tag_regs1_62;
      end else begin
        tag_regs1_56 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_57 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h39 == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_57 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_57 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_57 <= tag_regs1_62;
      end else begin
        tag_regs1_57 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_58 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h3a == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_58 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_58 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_58 <= tag_regs1_62;
      end else begin
        tag_regs1_58 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_59 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h3b == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_59 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_59 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_59 <= tag_regs1_62;
      end else begin
        tag_regs1_59 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_60 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h3c == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_60 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_60 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_60 <= tag_regs1_62;
      end else begin
        tag_regs1_60 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_61 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h3d == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_61 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_61 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[11:6]) begin
        tag_regs1_61 <= tag_regs1_62;
      end else begin
        tag_regs1_61 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_62 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h3e == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_62 <= io_wdata;
      end else if (6'h3f == io_waddr[11:6]) begin
        tag_regs1_62 <= tag_regs1_63;
      end else if (!(6'h3e == io_waddr[11:6])) begin
        tag_regs1_62 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 35:31]
      tag_regs1_63 <= 21'h0; // @[dcache_tag.scala 35:{37,37,37,37,37}]
    end else if (6'h3f == io_waddr[11:6]) begin // @[dcache_tag.scala 31:28]
      if (io_wen & io_waddr[5]) begin
        tag_regs1_63 <= io_wdata;
      end else if (!(6'h3f == io_waddr[11:6])) begin
        if (6'h3e == io_waddr[11:6]) begin
          tag_regs1_63 <= tag_regs1_62;
        end else begin
          tag_regs1_63 <= _GEN_189;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_regs0_0 = _RAND_0[20:0];
  _RAND_1 = {1{`RANDOM}};
  tag_regs0_1 = _RAND_1[20:0];
  _RAND_2 = {1{`RANDOM}};
  tag_regs0_2 = _RAND_2[20:0];
  _RAND_3 = {1{`RANDOM}};
  tag_regs0_3 = _RAND_3[20:0];
  _RAND_4 = {1{`RANDOM}};
  tag_regs0_4 = _RAND_4[20:0];
  _RAND_5 = {1{`RANDOM}};
  tag_regs0_5 = _RAND_5[20:0];
  _RAND_6 = {1{`RANDOM}};
  tag_regs0_6 = _RAND_6[20:0];
  _RAND_7 = {1{`RANDOM}};
  tag_regs0_7 = _RAND_7[20:0];
  _RAND_8 = {1{`RANDOM}};
  tag_regs0_8 = _RAND_8[20:0];
  _RAND_9 = {1{`RANDOM}};
  tag_regs0_9 = _RAND_9[20:0];
  _RAND_10 = {1{`RANDOM}};
  tag_regs0_10 = _RAND_10[20:0];
  _RAND_11 = {1{`RANDOM}};
  tag_regs0_11 = _RAND_11[20:0];
  _RAND_12 = {1{`RANDOM}};
  tag_regs0_12 = _RAND_12[20:0];
  _RAND_13 = {1{`RANDOM}};
  tag_regs0_13 = _RAND_13[20:0];
  _RAND_14 = {1{`RANDOM}};
  tag_regs0_14 = _RAND_14[20:0];
  _RAND_15 = {1{`RANDOM}};
  tag_regs0_15 = _RAND_15[20:0];
  _RAND_16 = {1{`RANDOM}};
  tag_regs0_16 = _RAND_16[20:0];
  _RAND_17 = {1{`RANDOM}};
  tag_regs0_17 = _RAND_17[20:0];
  _RAND_18 = {1{`RANDOM}};
  tag_regs0_18 = _RAND_18[20:0];
  _RAND_19 = {1{`RANDOM}};
  tag_regs0_19 = _RAND_19[20:0];
  _RAND_20 = {1{`RANDOM}};
  tag_regs0_20 = _RAND_20[20:0];
  _RAND_21 = {1{`RANDOM}};
  tag_regs0_21 = _RAND_21[20:0];
  _RAND_22 = {1{`RANDOM}};
  tag_regs0_22 = _RAND_22[20:0];
  _RAND_23 = {1{`RANDOM}};
  tag_regs0_23 = _RAND_23[20:0];
  _RAND_24 = {1{`RANDOM}};
  tag_regs0_24 = _RAND_24[20:0];
  _RAND_25 = {1{`RANDOM}};
  tag_regs0_25 = _RAND_25[20:0];
  _RAND_26 = {1{`RANDOM}};
  tag_regs0_26 = _RAND_26[20:0];
  _RAND_27 = {1{`RANDOM}};
  tag_regs0_27 = _RAND_27[20:0];
  _RAND_28 = {1{`RANDOM}};
  tag_regs0_28 = _RAND_28[20:0];
  _RAND_29 = {1{`RANDOM}};
  tag_regs0_29 = _RAND_29[20:0];
  _RAND_30 = {1{`RANDOM}};
  tag_regs0_30 = _RAND_30[20:0];
  _RAND_31 = {1{`RANDOM}};
  tag_regs0_31 = _RAND_31[20:0];
  _RAND_32 = {1{`RANDOM}};
  tag_regs0_32 = _RAND_32[20:0];
  _RAND_33 = {1{`RANDOM}};
  tag_regs0_33 = _RAND_33[20:0];
  _RAND_34 = {1{`RANDOM}};
  tag_regs0_34 = _RAND_34[20:0];
  _RAND_35 = {1{`RANDOM}};
  tag_regs0_35 = _RAND_35[20:0];
  _RAND_36 = {1{`RANDOM}};
  tag_regs0_36 = _RAND_36[20:0];
  _RAND_37 = {1{`RANDOM}};
  tag_regs0_37 = _RAND_37[20:0];
  _RAND_38 = {1{`RANDOM}};
  tag_regs0_38 = _RAND_38[20:0];
  _RAND_39 = {1{`RANDOM}};
  tag_regs0_39 = _RAND_39[20:0];
  _RAND_40 = {1{`RANDOM}};
  tag_regs0_40 = _RAND_40[20:0];
  _RAND_41 = {1{`RANDOM}};
  tag_regs0_41 = _RAND_41[20:0];
  _RAND_42 = {1{`RANDOM}};
  tag_regs0_42 = _RAND_42[20:0];
  _RAND_43 = {1{`RANDOM}};
  tag_regs0_43 = _RAND_43[20:0];
  _RAND_44 = {1{`RANDOM}};
  tag_regs0_44 = _RAND_44[20:0];
  _RAND_45 = {1{`RANDOM}};
  tag_regs0_45 = _RAND_45[20:0];
  _RAND_46 = {1{`RANDOM}};
  tag_regs0_46 = _RAND_46[20:0];
  _RAND_47 = {1{`RANDOM}};
  tag_regs0_47 = _RAND_47[20:0];
  _RAND_48 = {1{`RANDOM}};
  tag_regs0_48 = _RAND_48[20:0];
  _RAND_49 = {1{`RANDOM}};
  tag_regs0_49 = _RAND_49[20:0];
  _RAND_50 = {1{`RANDOM}};
  tag_regs0_50 = _RAND_50[20:0];
  _RAND_51 = {1{`RANDOM}};
  tag_regs0_51 = _RAND_51[20:0];
  _RAND_52 = {1{`RANDOM}};
  tag_regs0_52 = _RAND_52[20:0];
  _RAND_53 = {1{`RANDOM}};
  tag_regs0_53 = _RAND_53[20:0];
  _RAND_54 = {1{`RANDOM}};
  tag_regs0_54 = _RAND_54[20:0];
  _RAND_55 = {1{`RANDOM}};
  tag_regs0_55 = _RAND_55[20:0];
  _RAND_56 = {1{`RANDOM}};
  tag_regs0_56 = _RAND_56[20:0];
  _RAND_57 = {1{`RANDOM}};
  tag_regs0_57 = _RAND_57[20:0];
  _RAND_58 = {1{`RANDOM}};
  tag_regs0_58 = _RAND_58[20:0];
  _RAND_59 = {1{`RANDOM}};
  tag_regs0_59 = _RAND_59[20:0];
  _RAND_60 = {1{`RANDOM}};
  tag_regs0_60 = _RAND_60[20:0];
  _RAND_61 = {1{`RANDOM}};
  tag_regs0_61 = _RAND_61[20:0];
  _RAND_62 = {1{`RANDOM}};
  tag_regs0_62 = _RAND_62[20:0];
  _RAND_63 = {1{`RANDOM}};
  tag_regs0_63 = _RAND_63[20:0];
  _RAND_64 = {1{`RANDOM}};
  tag_regs1_0 = _RAND_64[20:0];
  _RAND_65 = {1{`RANDOM}};
  tag_regs1_1 = _RAND_65[20:0];
  _RAND_66 = {1{`RANDOM}};
  tag_regs1_2 = _RAND_66[20:0];
  _RAND_67 = {1{`RANDOM}};
  tag_regs1_3 = _RAND_67[20:0];
  _RAND_68 = {1{`RANDOM}};
  tag_regs1_4 = _RAND_68[20:0];
  _RAND_69 = {1{`RANDOM}};
  tag_regs1_5 = _RAND_69[20:0];
  _RAND_70 = {1{`RANDOM}};
  tag_regs1_6 = _RAND_70[20:0];
  _RAND_71 = {1{`RANDOM}};
  tag_regs1_7 = _RAND_71[20:0];
  _RAND_72 = {1{`RANDOM}};
  tag_regs1_8 = _RAND_72[20:0];
  _RAND_73 = {1{`RANDOM}};
  tag_regs1_9 = _RAND_73[20:0];
  _RAND_74 = {1{`RANDOM}};
  tag_regs1_10 = _RAND_74[20:0];
  _RAND_75 = {1{`RANDOM}};
  tag_regs1_11 = _RAND_75[20:0];
  _RAND_76 = {1{`RANDOM}};
  tag_regs1_12 = _RAND_76[20:0];
  _RAND_77 = {1{`RANDOM}};
  tag_regs1_13 = _RAND_77[20:0];
  _RAND_78 = {1{`RANDOM}};
  tag_regs1_14 = _RAND_78[20:0];
  _RAND_79 = {1{`RANDOM}};
  tag_regs1_15 = _RAND_79[20:0];
  _RAND_80 = {1{`RANDOM}};
  tag_regs1_16 = _RAND_80[20:0];
  _RAND_81 = {1{`RANDOM}};
  tag_regs1_17 = _RAND_81[20:0];
  _RAND_82 = {1{`RANDOM}};
  tag_regs1_18 = _RAND_82[20:0];
  _RAND_83 = {1{`RANDOM}};
  tag_regs1_19 = _RAND_83[20:0];
  _RAND_84 = {1{`RANDOM}};
  tag_regs1_20 = _RAND_84[20:0];
  _RAND_85 = {1{`RANDOM}};
  tag_regs1_21 = _RAND_85[20:0];
  _RAND_86 = {1{`RANDOM}};
  tag_regs1_22 = _RAND_86[20:0];
  _RAND_87 = {1{`RANDOM}};
  tag_regs1_23 = _RAND_87[20:0];
  _RAND_88 = {1{`RANDOM}};
  tag_regs1_24 = _RAND_88[20:0];
  _RAND_89 = {1{`RANDOM}};
  tag_regs1_25 = _RAND_89[20:0];
  _RAND_90 = {1{`RANDOM}};
  tag_regs1_26 = _RAND_90[20:0];
  _RAND_91 = {1{`RANDOM}};
  tag_regs1_27 = _RAND_91[20:0];
  _RAND_92 = {1{`RANDOM}};
  tag_regs1_28 = _RAND_92[20:0];
  _RAND_93 = {1{`RANDOM}};
  tag_regs1_29 = _RAND_93[20:0];
  _RAND_94 = {1{`RANDOM}};
  tag_regs1_30 = _RAND_94[20:0];
  _RAND_95 = {1{`RANDOM}};
  tag_regs1_31 = _RAND_95[20:0];
  _RAND_96 = {1{`RANDOM}};
  tag_regs1_32 = _RAND_96[20:0];
  _RAND_97 = {1{`RANDOM}};
  tag_regs1_33 = _RAND_97[20:0];
  _RAND_98 = {1{`RANDOM}};
  tag_regs1_34 = _RAND_98[20:0];
  _RAND_99 = {1{`RANDOM}};
  tag_regs1_35 = _RAND_99[20:0];
  _RAND_100 = {1{`RANDOM}};
  tag_regs1_36 = _RAND_100[20:0];
  _RAND_101 = {1{`RANDOM}};
  tag_regs1_37 = _RAND_101[20:0];
  _RAND_102 = {1{`RANDOM}};
  tag_regs1_38 = _RAND_102[20:0];
  _RAND_103 = {1{`RANDOM}};
  tag_regs1_39 = _RAND_103[20:0];
  _RAND_104 = {1{`RANDOM}};
  tag_regs1_40 = _RAND_104[20:0];
  _RAND_105 = {1{`RANDOM}};
  tag_regs1_41 = _RAND_105[20:0];
  _RAND_106 = {1{`RANDOM}};
  tag_regs1_42 = _RAND_106[20:0];
  _RAND_107 = {1{`RANDOM}};
  tag_regs1_43 = _RAND_107[20:0];
  _RAND_108 = {1{`RANDOM}};
  tag_regs1_44 = _RAND_108[20:0];
  _RAND_109 = {1{`RANDOM}};
  tag_regs1_45 = _RAND_109[20:0];
  _RAND_110 = {1{`RANDOM}};
  tag_regs1_46 = _RAND_110[20:0];
  _RAND_111 = {1{`RANDOM}};
  tag_regs1_47 = _RAND_111[20:0];
  _RAND_112 = {1{`RANDOM}};
  tag_regs1_48 = _RAND_112[20:0];
  _RAND_113 = {1{`RANDOM}};
  tag_regs1_49 = _RAND_113[20:0];
  _RAND_114 = {1{`RANDOM}};
  tag_regs1_50 = _RAND_114[20:0];
  _RAND_115 = {1{`RANDOM}};
  tag_regs1_51 = _RAND_115[20:0];
  _RAND_116 = {1{`RANDOM}};
  tag_regs1_52 = _RAND_116[20:0];
  _RAND_117 = {1{`RANDOM}};
  tag_regs1_53 = _RAND_117[20:0];
  _RAND_118 = {1{`RANDOM}};
  tag_regs1_54 = _RAND_118[20:0];
  _RAND_119 = {1{`RANDOM}};
  tag_regs1_55 = _RAND_119[20:0];
  _RAND_120 = {1{`RANDOM}};
  tag_regs1_56 = _RAND_120[20:0];
  _RAND_121 = {1{`RANDOM}};
  tag_regs1_57 = _RAND_121[20:0];
  _RAND_122 = {1{`RANDOM}};
  tag_regs1_58 = _RAND_122[20:0];
  _RAND_123 = {1{`RANDOM}};
  tag_regs1_59 = _RAND_123[20:0];
  _RAND_124 = {1{`RANDOM}};
  tag_regs1_60 = _RAND_124[20:0];
  _RAND_125 = {1{`RANDOM}};
  tag_regs1_61 = _RAND_125[20:0];
  _RAND_126 = {1{`RANDOM}};
  tag_regs1_62 = _RAND_126[20:0];
  _RAND_127 = {1{`RANDOM}};
  tag_regs1_63 = _RAND_127[20:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    tag_regs0_0 = 21'h0;
  end
  if (reset) begin
    tag_regs0_1 = 21'h0;
  end
  if (reset) begin
    tag_regs0_2 = 21'h0;
  end
  if (reset) begin
    tag_regs0_3 = 21'h0;
  end
  if (reset) begin
    tag_regs0_4 = 21'h0;
  end
  if (reset) begin
    tag_regs0_5 = 21'h0;
  end
  if (reset) begin
    tag_regs0_6 = 21'h0;
  end
  if (reset) begin
    tag_regs0_7 = 21'h0;
  end
  if (reset) begin
    tag_regs0_8 = 21'h0;
  end
  if (reset) begin
    tag_regs0_9 = 21'h0;
  end
  if (reset) begin
    tag_regs0_10 = 21'h0;
  end
  if (reset) begin
    tag_regs0_11 = 21'h0;
  end
  if (reset) begin
    tag_regs0_12 = 21'h0;
  end
  if (reset) begin
    tag_regs0_13 = 21'h0;
  end
  if (reset) begin
    tag_regs0_14 = 21'h0;
  end
  if (reset) begin
    tag_regs0_15 = 21'h0;
  end
  if (reset) begin
    tag_regs0_16 = 21'h0;
  end
  if (reset) begin
    tag_regs0_17 = 21'h0;
  end
  if (reset) begin
    tag_regs0_18 = 21'h0;
  end
  if (reset) begin
    tag_regs0_19 = 21'h0;
  end
  if (reset) begin
    tag_regs0_20 = 21'h0;
  end
  if (reset) begin
    tag_regs0_21 = 21'h0;
  end
  if (reset) begin
    tag_regs0_22 = 21'h0;
  end
  if (reset) begin
    tag_regs0_23 = 21'h0;
  end
  if (reset) begin
    tag_regs0_24 = 21'h0;
  end
  if (reset) begin
    tag_regs0_25 = 21'h0;
  end
  if (reset) begin
    tag_regs0_26 = 21'h0;
  end
  if (reset) begin
    tag_regs0_27 = 21'h0;
  end
  if (reset) begin
    tag_regs0_28 = 21'h0;
  end
  if (reset) begin
    tag_regs0_29 = 21'h0;
  end
  if (reset) begin
    tag_regs0_30 = 21'h0;
  end
  if (reset) begin
    tag_regs0_31 = 21'h0;
  end
  if (reset) begin
    tag_regs0_32 = 21'h0;
  end
  if (reset) begin
    tag_regs0_33 = 21'h0;
  end
  if (reset) begin
    tag_regs0_34 = 21'h0;
  end
  if (reset) begin
    tag_regs0_35 = 21'h0;
  end
  if (reset) begin
    tag_regs0_36 = 21'h0;
  end
  if (reset) begin
    tag_regs0_37 = 21'h0;
  end
  if (reset) begin
    tag_regs0_38 = 21'h0;
  end
  if (reset) begin
    tag_regs0_39 = 21'h0;
  end
  if (reset) begin
    tag_regs0_40 = 21'h0;
  end
  if (reset) begin
    tag_regs0_41 = 21'h0;
  end
  if (reset) begin
    tag_regs0_42 = 21'h0;
  end
  if (reset) begin
    tag_regs0_43 = 21'h0;
  end
  if (reset) begin
    tag_regs0_44 = 21'h0;
  end
  if (reset) begin
    tag_regs0_45 = 21'h0;
  end
  if (reset) begin
    tag_regs0_46 = 21'h0;
  end
  if (reset) begin
    tag_regs0_47 = 21'h0;
  end
  if (reset) begin
    tag_regs0_48 = 21'h0;
  end
  if (reset) begin
    tag_regs0_49 = 21'h0;
  end
  if (reset) begin
    tag_regs0_50 = 21'h0;
  end
  if (reset) begin
    tag_regs0_51 = 21'h0;
  end
  if (reset) begin
    tag_regs0_52 = 21'h0;
  end
  if (reset) begin
    tag_regs0_53 = 21'h0;
  end
  if (reset) begin
    tag_regs0_54 = 21'h0;
  end
  if (reset) begin
    tag_regs0_55 = 21'h0;
  end
  if (reset) begin
    tag_regs0_56 = 21'h0;
  end
  if (reset) begin
    tag_regs0_57 = 21'h0;
  end
  if (reset) begin
    tag_regs0_58 = 21'h0;
  end
  if (reset) begin
    tag_regs0_59 = 21'h0;
  end
  if (reset) begin
    tag_regs0_60 = 21'h0;
  end
  if (reset) begin
    tag_regs0_61 = 21'h0;
  end
  if (reset) begin
    tag_regs0_62 = 21'h0;
  end
  if (reset) begin
    tag_regs0_63 = 21'h0;
  end
  if (reset) begin
    tag_regs1_0 = 21'h0;
  end
  if (reset) begin
    tag_regs1_1 = 21'h0;
  end
  if (reset) begin
    tag_regs1_2 = 21'h0;
  end
  if (reset) begin
    tag_regs1_3 = 21'h0;
  end
  if (reset) begin
    tag_regs1_4 = 21'h0;
  end
  if (reset) begin
    tag_regs1_5 = 21'h0;
  end
  if (reset) begin
    tag_regs1_6 = 21'h0;
  end
  if (reset) begin
    tag_regs1_7 = 21'h0;
  end
  if (reset) begin
    tag_regs1_8 = 21'h0;
  end
  if (reset) begin
    tag_regs1_9 = 21'h0;
  end
  if (reset) begin
    tag_regs1_10 = 21'h0;
  end
  if (reset) begin
    tag_regs1_11 = 21'h0;
  end
  if (reset) begin
    tag_regs1_12 = 21'h0;
  end
  if (reset) begin
    tag_regs1_13 = 21'h0;
  end
  if (reset) begin
    tag_regs1_14 = 21'h0;
  end
  if (reset) begin
    tag_regs1_15 = 21'h0;
  end
  if (reset) begin
    tag_regs1_16 = 21'h0;
  end
  if (reset) begin
    tag_regs1_17 = 21'h0;
  end
  if (reset) begin
    tag_regs1_18 = 21'h0;
  end
  if (reset) begin
    tag_regs1_19 = 21'h0;
  end
  if (reset) begin
    tag_regs1_20 = 21'h0;
  end
  if (reset) begin
    tag_regs1_21 = 21'h0;
  end
  if (reset) begin
    tag_regs1_22 = 21'h0;
  end
  if (reset) begin
    tag_regs1_23 = 21'h0;
  end
  if (reset) begin
    tag_regs1_24 = 21'h0;
  end
  if (reset) begin
    tag_regs1_25 = 21'h0;
  end
  if (reset) begin
    tag_regs1_26 = 21'h0;
  end
  if (reset) begin
    tag_regs1_27 = 21'h0;
  end
  if (reset) begin
    tag_regs1_28 = 21'h0;
  end
  if (reset) begin
    tag_regs1_29 = 21'h0;
  end
  if (reset) begin
    tag_regs1_30 = 21'h0;
  end
  if (reset) begin
    tag_regs1_31 = 21'h0;
  end
  if (reset) begin
    tag_regs1_32 = 21'h0;
  end
  if (reset) begin
    tag_regs1_33 = 21'h0;
  end
  if (reset) begin
    tag_regs1_34 = 21'h0;
  end
  if (reset) begin
    tag_regs1_35 = 21'h0;
  end
  if (reset) begin
    tag_regs1_36 = 21'h0;
  end
  if (reset) begin
    tag_regs1_37 = 21'h0;
  end
  if (reset) begin
    tag_regs1_38 = 21'h0;
  end
  if (reset) begin
    tag_regs1_39 = 21'h0;
  end
  if (reset) begin
    tag_regs1_40 = 21'h0;
  end
  if (reset) begin
    tag_regs1_41 = 21'h0;
  end
  if (reset) begin
    tag_regs1_42 = 21'h0;
  end
  if (reset) begin
    tag_regs1_43 = 21'h0;
  end
  if (reset) begin
    tag_regs1_44 = 21'h0;
  end
  if (reset) begin
    tag_regs1_45 = 21'h0;
  end
  if (reset) begin
    tag_regs1_46 = 21'h0;
  end
  if (reset) begin
    tag_regs1_47 = 21'h0;
  end
  if (reset) begin
    tag_regs1_48 = 21'h0;
  end
  if (reset) begin
    tag_regs1_49 = 21'h0;
  end
  if (reset) begin
    tag_regs1_50 = 21'h0;
  end
  if (reset) begin
    tag_regs1_51 = 21'h0;
  end
  if (reset) begin
    tag_regs1_52 = 21'h0;
  end
  if (reset) begin
    tag_regs1_53 = 21'h0;
  end
  if (reset) begin
    tag_regs1_54 = 21'h0;
  end
  if (reset) begin
    tag_regs1_55 = 21'h0;
  end
  if (reset) begin
    tag_regs1_56 = 21'h0;
  end
  if (reset) begin
    tag_regs1_57 = 21'h0;
  end
  if (reset) begin
    tag_regs1_58 = 21'h0;
  end
  if (reset) begin
    tag_regs1_59 = 21'h0;
  end
  if (reset) begin
    tag_regs1_60 = 21'h0;
  end
  if (reset) begin
    tag_regs1_61 = 21'h0;
  end
  if (reset) begin
    tag_regs1_62 = 21'h0;
  end
  if (reset) begin
    tag_regs1_63 = 21'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module dcache_data(
  input         clock,
  input  [3:0]  io_wen,
  input  [31:0] io_addr,
  input  [31:0] io_wdata,
  output [31:0] io_rdata
);
  wire  dcache_data_ram_0_clka; // @[dcache_data.scala 32:35]
  wire  dcache_data_ram_0_ena; // @[dcache_data.scala 32:35]
  wire [3:0] dcache_data_ram_0_wea; // @[dcache_data.scala 32:35]
  wire [6:0] dcache_data_ram_0_addra; // @[dcache_data.scala 32:35]
  wire [31:0] dcache_data_ram_0_dina; // @[dcache_data.scala 32:35]
  wire [31:0] dcache_data_ram_0_douta; // @[dcache_data.scala 32:35]
  dcache_data_ram dcache_data_ram_0 ( // @[dcache_data.scala 32:35]
    .clka(dcache_data_ram_0_clka),
    .ena(dcache_data_ram_0_ena),
    .wea(dcache_data_ram_0_wea),
    .addra(dcache_data_ram_0_addra),
    .dina(dcache_data_ram_0_dina),
    .douta(dcache_data_ram_0_douta)
  );
  assign io_rdata = dcache_data_ram_0_douta; // @[dcache_data.scala 38:18]
  assign dcache_data_ram_0_clka = clock; // @[dcache_data.scala 33:40]
  assign dcache_data_ram_0_ena = 1'h1; // @[dcache_data.scala 34:32]
  assign dcache_data_ram_0_wea = io_wen; // @[dcache_data.scala 35:31]
  assign dcache_data_ram_0_addra = io_addr[11:5]; // @[dcache_data.scala 36:42]
  assign dcache_data_ram_0_dina = io_wdata; // @[dcache_data.scala 37:31]
endmodule
module data_cache(
  input         clock,
  input         reset,
  output [31:0] io_port_araddr,
  output [3:0]  io_port_arlen,
  output [2:0]  io_port_arsize,
  output [1:0]  io_port_arburst,
  output        io_port_arvalid,
  input         io_port_arready,
  input  [31:0] io_port_rdata,
  input         io_port_rlast,
  input         io_port_rvalid,
  output [31:0] io_port_awaddr,
  output [3:0]  io_port_awlen,
  output [2:0]  io_port_awsize,
  output [1:0]  io_port_awburst,
  output        io_port_awvalid,
  input         io_port_awready,
  output [31:0] io_port_wdata,
  output [3:0]  io_port_wstrb,
  output        io_port_wlast,
  output        io_port_wvalid,
  input         io_port_wready,
  input         io_port_bvalid,
  input         io_port_sram_req,
  input         io_port_sram_wr,
  input  [1:0]  io_port_sram_size,
  input  [31:0] io_port_sram_addr,
  input  [31:0] io_port_sram_wdata,
  output [31:0] io_port_sram_rdata,
  input         io_port_sram_cache,
  output        io_stage2_stall,
  output        io_stage1_wr,
  output [31:0] io_v_addr_for_tlb,
  input  [31:0] io_p_addr_for_tlb,
  output        io_tlb_req,
  input  [2:0]  io_tlb_exception,
  output [2:0]  io_stage1_tlb_exception,
  input  [3:0]  io_data_wstrb
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
`endif // RANDOMIZE_REG_INIT
  wire  dcache_tag_clock; // @[data_cache.scala 37:30]
  wire  dcache_tag_reset; // @[data_cache.scala 37:30]
  wire  dcache_tag_io_wen; // @[data_cache.scala 37:30]
  wire [20:0] dcache_tag_io_wdata; // @[data_cache.scala 37:30]
  wire [31:0] dcache_tag_io_raddr; // @[data_cache.scala 37:30]
  wire [31:0] dcache_tag_io_waddr; // @[data_cache.scala 37:30]
  wire  dcache_tag_io_hit; // @[data_cache.scala 37:30]
  wire  dcache_tag_io_valid; // @[data_cache.scala 37:30]
  wire [19:0] dcache_tag_io_tag; // @[data_cache.scala 37:30]
  wire  dcache_tag_1_clock; // @[data_cache.scala 38:30]
  wire  dcache_tag_1_reset; // @[data_cache.scala 38:30]
  wire  dcache_tag_1_io_wen; // @[data_cache.scala 38:30]
  wire [20:0] dcache_tag_1_io_wdata; // @[data_cache.scala 38:30]
  wire [31:0] dcache_tag_1_io_raddr; // @[data_cache.scala 38:30]
  wire [31:0] dcache_tag_1_io_waddr; // @[data_cache.scala 38:30]
  wire  dcache_tag_1_io_hit; // @[data_cache.scala 38:30]
  wire  dcache_tag_1_io_valid; // @[data_cache.scala 38:30]
  wire [19:0] dcache_tag_1_io_tag; // @[data_cache.scala 38:30]
  wire  dcache_data_clock; // @[data_cache.scala 70:55]
  wire [3:0] dcache_data_io_wen; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_io_addr; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_io_wdata; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_io_rdata; // @[data_cache.scala 70:55]
  wire  dcache_data_1_clock; // @[data_cache.scala 70:55]
  wire [3:0] dcache_data_1_io_wen; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_1_io_addr; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_1_io_wdata; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_1_io_rdata; // @[data_cache.scala 70:55]
  wire  dcache_data_2_clock; // @[data_cache.scala 70:55]
  wire [3:0] dcache_data_2_io_wen; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_2_io_addr; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_2_io_wdata; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_2_io_rdata; // @[data_cache.scala 70:55]
  wire  dcache_data_3_clock; // @[data_cache.scala 70:55]
  wire [3:0] dcache_data_3_io_wen; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_3_io_addr; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_3_io_wdata; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_3_io_rdata; // @[data_cache.scala 70:55]
  wire  dcache_data_4_clock; // @[data_cache.scala 70:55]
  wire [3:0] dcache_data_4_io_wen; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_4_io_addr; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_4_io_wdata; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_4_io_rdata; // @[data_cache.scala 70:55]
  wire  dcache_data_5_clock; // @[data_cache.scala 70:55]
  wire [3:0] dcache_data_5_io_wen; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_5_io_addr; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_5_io_wdata; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_5_io_rdata; // @[data_cache.scala 70:55]
  wire  dcache_data_6_clock; // @[data_cache.scala 70:55]
  wire [3:0] dcache_data_6_io_wen; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_6_io_addr; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_6_io_wdata; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_6_io_rdata; // @[data_cache.scala 70:55]
  wire  dcache_data_7_clock; // @[data_cache.scala 70:55]
  wire [3:0] dcache_data_7_io_wen; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_7_io_addr; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_7_io_wdata; // @[data_cache.scala 70:55]
  wire [31:0] dcache_data_7_io_rdata; // @[data_cache.scala 70:55]
  wire  dcache_data_8_clock; // @[data_cache.scala 71:55]
  wire [3:0] dcache_data_8_io_wen; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_8_io_addr; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_8_io_wdata; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_8_io_rdata; // @[data_cache.scala 71:55]
  wire  dcache_data_9_clock; // @[data_cache.scala 71:55]
  wire [3:0] dcache_data_9_io_wen; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_9_io_addr; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_9_io_wdata; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_9_io_rdata; // @[data_cache.scala 71:55]
  wire  dcache_data_10_clock; // @[data_cache.scala 71:55]
  wire [3:0] dcache_data_10_io_wen; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_10_io_addr; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_10_io_wdata; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_10_io_rdata; // @[data_cache.scala 71:55]
  wire  dcache_data_11_clock; // @[data_cache.scala 71:55]
  wire [3:0] dcache_data_11_io_wen; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_11_io_addr; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_11_io_wdata; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_11_io_rdata; // @[data_cache.scala 71:55]
  wire  dcache_data_12_clock; // @[data_cache.scala 71:55]
  wire [3:0] dcache_data_12_io_wen; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_12_io_addr; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_12_io_wdata; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_12_io_rdata; // @[data_cache.scala 71:55]
  wire  dcache_data_13_clock; // @[data_cache.scala 71:55]
  wire [3:0] dcache_data_13_io_wen; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_13_io_addr; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_13_io_wdata; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_13_io_rdata; // @[data_cache.scala 71:55]
  wire  dcache_data_14_clock; // @[data_cache.scala 71:55]
  wire [3:0] dcache_data_14_io_wen; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_14_io_addr; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_14_io_wdata; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_14_io_rdata; // @[data_cache.scala 71:55]
  wire  dcache_data_15_clock; // @[data_cache.scala 71:55]
  wire [3:0] dcache_data_15_io_wen; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_15_io_addr; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_15_io_wdata; // @[data_cache.scala 71:55]
  wire [31:0] dcache_data_15_io_rdata; // @[data_cache.scala 71:55]
  reg [4:0] work_state; // @[data_cache.scala 30:29]
  reg [2:0] write_counter; // @[data_cache.scala 32:33]
  reg [2:0] read_counter; // @[data_cache.scala 33:32]
  reg [31:0] wait_data; // @[data_cache.scala 34:29]
  reg  lru_0; // @[data_cache.scala 40:22]
  reg  lru_1; // @[data_cache.scala 40:22]
  reg  lru_2; // @[data_cache.scala 40:22]
  reg  lru_3; // @[data_cache.scala 40:22]
  reg  lru_4; // @[data_cache.scala 40:22]
  reg  lru_5; // @[data_cache.scala 40:22]
  reg  lru_6; // @[data_cache.scala 40:22]
  reg  lru_7; // @[data_cache.scala 40:22]
  reg  lru_8; // @[data_cache.scala 40:22]
  reg  lru_9; // @[data_cache.scala 40:22]
  reg  lru_10; // @[data_cache.scala 40:22]
  reg  lru_11; // @[data_cache.scala 40:22]
  reg  lru_12; // @[data_cache.scala 40:22]
  reg  lru_13; // @[data_cache.scala 40:22]
  reg  lru_14; // @[data_cache.scala 40:22]
  reg  lru_15; // @[data_cache.scala 40:22]
  reg  lru_16; // @[data_cache.scala 40:22]
  reg  lru_17; // @[data_cache.scala 40:22]
  reg  lru_18; // @[data_cache.scala 40:22]
  reg  lru_19; // @[data_cache.scala 40:22]
  reg  lru_20; // @[data_cache.scala 40:22]
  reg  lru_21; // @[data_cache.scala 40:22]
  reg  lru_22; // @[data_cache.scala 40:22]
  reg  lru_23; // @[data_cache.scala 40:22]
  reg  lru_24; // @[data_cache.scala 40:22]
  reg  lru_25; // @[data_cache.scala 40:22]
  reg  lru_26; // @[data_cache.scala 40:22]
  reg  lru_27; // @[data_cache.scala 40:22]
  reg  lru_28; // @[data_cache.scala 40:22]
  reg  lru_29; // @[data_cache.scala 40:22]
  reg  lru_30; // @[data_cache.scala 40:22]
  reg  lru_31; // @[data_cache.scala 40:22]
  reg  lru_32; // @[data_cache.scala 40:22]
  reg  lru_33; // @[data_cache.scala 40:22]
  reg  lru_34; // @[data_cache.scala 40:22]
  reg  lru_35; // @[data_cache.scala 40:22]
  reg  lru_36; // @[data_cache.scala 40:22]
  reg  lru_37; // @[data_cache.scala 40:22]
  reg  lru_38; // @[data_cache.scala 40:22]
  reg  lru_39; // @[data_cache.scala 40:22]
  reg  lru_40; // @[data_cache.scala 40:22]
  reg  lru_41; // @[data_cache.scala 40:22]
  reg  lru_42; // @[data_cache.scala 40:22]
  reg  lru_43; // @[data_cache.scala 40:22]
  reg  lru_44; // @[data_cache.scala 40:22]
  reg  lru_45; // @[data_cache.scala 40:22]
  reg  lru_46; // @[data_cache.scala 40:22]
  reg  lru_47; // @[data_cache.scala 40:22]
  reg  lru_48; // @[data_cache.scala 40:22]
  reg  lru_49; // @[data_cache.scala 40:22]
  reg  lru_50; // @[data_cache.scala 40:22]
  reg  lru_51; // @[data_cache.scala 40:22]
  reg  lru_52; // @[data_cache.scala 40:22]
  reg  lru_53; // @[data_cache.scala 40:22]
  reg  lru_54; // @[data_cache.scala 40:22]
  reg  lru_55; // @[data_cache.scala 40:22]
  reg  lru_56; // @[data_cache.scala 40:22]
  reg  lru_57; // @[data_cache.scala 40:22]
  reg  lru_58; // @[data_cache.scala 40:22]
  reg  lru_59; // @[data_cache.scala 40:22]
  reg  lru_60; // @[data_cache.scala 40:22]
  reg  lru_61; // @[data_cache.scala 40:22]
  reg  lru_62; // @[data_cache.scala 40:22]
  reg  lru_63; // @[data_cache.scala 40:22]
  reg  lru_64; // @[data_cache.scala 40:22]
  reg  lru_65; // @[data_cache.scala 40:22]
  reg  lru_66; // @[data_cache.scala 40:22]
  reg  lru_67; // @[data_cache.scala 40:22]
  reg  lru_68; // @[data_cache.scala 40:22]
  reg  lru_69; // @[data_cache.scala 40:22]
  reg  lru_70; // @[data_cache.scala 40:22]
  reg  lru_71; // @[data_cache.scala 40:22]
  reg  lru_72; // @[data_cache.scala 40:22]
  reg  lru_73; // @[data_cache.scala 40:22]
  reg  lru_74; // @[data_cache.scala 40:22]
  reg  lru_75; // @[data_cache.scala 40:22]
  reg  lru_76; // @[data_cache.scala 40:22]
  reg  lru_77; // @[data_cache.scala 40:22]
  reg  lru_78; // @[data_cache.scala 40:22]
  reg  lru_79; // @[data_cache.scala 40:22]
  reg  lru_80; // @[data_cache.scala 40:22]
  reg  lru_81; // @[data_cache.scala 40:22]
  reg  lru_82; // @[data_cache.scala 40:22]
  reg  lru_83; // @[data_cache.scala 40:22]
  reg  lru_84; // @[data_cache.scala 40:22]
  reg  lru_85; // @[data_cache.scala 40:22]
  reg  lru_86; // @[data_cache.scala 40:22]
  reg  lru_87; // @[data_cache.scala 40:22]
  reg  lru_88; // @[data_cache.scala 40:22]
  reg  lru_89; // @[data_cache.scala 40:22]
  reg  lru_90; // @[data_cache.scala 40:22]
  reg  lru_91; // @[data_cache.scala 40:22]
  reg  lru_92; // @[data_cache.scala 40:22]
  reg  lru_93; // @[data_cache.scala 40:22]
  reg  lru_94; // @[data_cache.scala 40:22]
  reg  lru_95; // @[data_cache.scala 40:22]
  reg  lru_96; // @[data_cache.scala 40:22]
  reg  lru_97; // @[data_cache.scala 40:22]
  reg  lru_98; // @[data_cache.scala 40:22]
  reg  lru_99; // @[data_cache.scala 40:22]
  reg  lru_100; // @[data_cache.scala 40:22]
  reg  lru_101; // @[data_cache.scala 40:22]
  reg  lru_102; // @[data_cache.scala 40:22]
  reg  lru_103; // @[data_cache.scala 40:22]
  reg  lru_104; // @[data_cache.scala 40:22]
  reg  lru_105; // @[data_cache.scala 40:22]
  reg  lru_106; // @[data_cache.scala 40:22]
  reg  lru_107; // @[data_cache.scala 40:22]
  reg  lru_108; // @[data_cache.scala 40:22]
  reg  lru_109; // @[data_cache.scala 40:22]
  reg  lru_110; // @[data_cache.scala 40:22]
  reg  lru_111; // @[data_cache.scala 40:22]
  reg  lru_112; // @[data_cache.scala 40:22]
  reg  lru_113; // @[data_cache.scala 40:22]
  reg  lru_114; // @[data_cache.scala 40:22]
  reg  lru_115; // @[data_cache.scala 40:22]
  reg  lru_116; // @[data_cache.scala 40:22]
  reg  lru_117; // @[data_cache.scala 40:22]
  reg  lru_118; // @[data_cache.scala 40:22]
  reg  lru_119; // @[data_cache.scala 40:22]
  reg  lru_120; // @[data_cache.scala 40:22]
  reg  lru_121; // @[data_cache.scala 40:22]
  reg  lru_122; // @[data_cache.scala 40:22]
  reg  lru_123; // @[data_cache.scala 40:22]
  reg  lru_124; // @[data_cache.scala 40:22]
  reg  lru_125; // @[data_cache.scala 40:22]
  reg  lru_126; // @[data_cache.scala 40:22]
  reg  lru_127; // @[data_cache.scala 40:22]
  reg  way0_dirty_0; // @[data_cache.scala 41:29]
  reg  way0_dirty_1; // @[data_cache.scala 41:29]
  reg  way0_dirty_2; // @[data_cache.scala 41:29]
  reg  way0_dirty_3; // @[data_cache.scala 41:29]
  reg  way0_dirty_4; // @[data_cache.scala 41:29]
  reg  way0_dirty_5; // @[data_cache.scala 41:29]
  reg  way0_dirty_6; // @[data_cache.scala 41:29]
  reg  way0_dirty_7; // @[data_cache.scala 41:29]
  reg  way0_dirty_8; // @[data_cache.scala 41:29]
  reg  way0_dirty_9; // @[data_cache.scala 41:29]
  reg  way0_dirty_10; // @[data_cache.scala 41:29]
  reg  way0_dirty_11; // @[data_cache.scala 41:29]
  reg  way0_dirty_12; // @[data_cache.scala 41:29]
  reg  way0_dirty_13; // @[data_cache.scala 41:29]
  reg  way0_dirty_14; // @[data_cache.scala 41:29]
  reg  way0_dirty_15; // @[data_cache.scala 41:29]
  reg  way0_dirty_16; // @[data_cache.scala 41:29]
  reg  way0_dirty_17; // @[data_cache.scala 41:29]
  reg  way0_dirty_18; // @[data_cache.scala 41:29]
  reg  way0_dirty_19; // @[data_cache.scala 41:29]
  reg  way0_dirty_20; // @[data_cache.scala 41:29]
  reg  way0_dirty_21; // @[data_cache.scala 41:29]
  reg  way0_dirty_22; // @[data_cache.scala 41:29]
  reg  way0_dirty_23; // @[data_cache.scala 41:29]
  reg  way0_dirty_24; // @[data_cache.scala 41:29]
  reg  way0_dirty_25; // @[data_cache.scala 41:29]
  reg  way0_dirty_26; // @[data_cache.scala 41:29]
  reg  way0_dirty_27; // @[data_cache.scala 41:29]
  reg  way0_dirty_28; // @[data_cache.scala 41:29]
  reg  way0_dirty_29; // @[data_cache.scala 41:29]
  reg  way0_dirty_30; // @[data_cache.scala 41:29]
  reg  way0_dirty_31; // @[data_cache.scala 41:29]
  reg  way0_dirty_32; // @[data_cache.scala 41:29]
  reg  way0_dirty_33; // @[data_cache.scala 41:29]
  reg  way0_dirty_34; // @[data_cache.scala 41:29]
  reg  way0_dirty_35; // @[data_cache.scala 41:29]
  reg  way0_dirty_36; // @[data_cache.scala 41:29]
  reg  way0_dirty_37; // @[data_cache.scala 41:29]
  reg  way0_dirty_38; // @[data_cache.scala 41:29]
  reg  way0_dirty_39; // @[data_cache.scala 41:29]
  reg  way0_dirty_40; // @[data_cache.scala 41:29]
  reg  way0_dirty_41; // @[data_cache.scala 41:29]
  reg  way0_dirty_42; // @[data_cache.scala 41:29]
  reg  way0_dirty_43; // @[data_cache.scala 41:29]
  reg  way0_dirty_44; // @[data_cache.scala 41:29]
  reg  way0_dirty_45; // @[data_cache.scala 41:29]
  reg  way0_dirty_46; // @[data_cache.scala 41:29]
  reg  way0_dirty_47; // @[data_cache.scala 41:29]
  reg  way0_dirty_48; // @[data_cache.scala 41:29]
  reg  way0_dirty_49; // @[data_cache.scala 41:29]
  reg  way0_dirty_50; // @[data_cache.scala 41:29]
  reg  way0_dirty_51; // @[data_cache.scala 41:29]
  reg  way0_dirty_52; // @[data_cache.scala 41:29]
  reg  way0_dirty_53; // @[data_cache.scala 41:29]
  reg  way0_dirty_54; // @[data_cache.scala 41:29]
  reg  way0_dirty_55; // @[data_cache.scala 41:29]
  reg  way0_dirty_56; // @[data_cache.scala 41:29]
  reg  way0_dirty_57; // @[data_cache.scala 41:29]
  reg  way0_dirty_58; // @[data_cache.scala 41:29]
  reg  way0_dirty_59; // @[data_cache.scala 41:29]
  reg  way0_dirty_60; // @[data_cache.scala 41:29]
  reg  way0_dirty_61; // @[data_cache.scala 41:29]
  reg  way0_dirty_62; // @[data_cache.scala 41:29]
  reg  way0_dirty_63; // @[data_cache.scala 41:29]
  reg  way0_dirty_64; // @[data_cache.scala 41:29]
  reg  way0_dirty_65; // @[data_cache.scala 41:29]
  reg  way0_dirty_66; // @[data_cache.scala 41:29]
  reg  way0_dirty_67; // @[data_cache.scala 41:29]
  reg  way0_dirty_68; // @[data_cache.scala 41:29]
  reg  way0_dirty_69; // @[data_cache.scala 41:29]
  reg  way0_dirty_70; // @[data_cache.scala 41:29]
  reg  way0_dirty_71; // @[data_cache.scala 41:29]
  reg  way0_dirty_72; // @[data_cache.scala 41:29]
  reg  way0_dirty_73; // @[data_cache.scala 41:29]
  reg  way0_dirty_74; // @[data_cache.scala 41:29]
  reg  way0_dirty_75; // @[data_cache.scala 41:29]
  reg  way0_dirty_76; // @[data_cache.scala 41:29]
  reg  way0_dirty_77; // @[data_cache.scala 41:29]
  reg  way0_dirty_78; // @[data_cache.scala 41:29]
  reg  way0_dirty_79; // @[data_cache.scala 41:29]
  reg  way0_dirty_80; // @[data_cache.scala 41:29]
  reg  way0_dirty_81; // @[data_cache.scala 41:29]
  reg  way0_dirty_82; // @[data_cache.scala 41:29]
  reg  way0_dirty_83; // @[data_cache.scala 41:29]
  reg  way0_dirty_84; // @[data_cache.scala 41:29]
  reg  way0_dirty_85; // @[data_cache.scala 41:29]
  reg  way0_dirty_86; // @[data_cache.scala 41:29]
  reg  way0_dirty_87; // @[data_cache.scala 41:29]
  reg  way0_dirty_88; // @[data_cache.scala 41:29]
  reg  way0_dirty_89; // @[data_cache.scala 41:29]
  reg  way0_dirty_90; // @[data_cache.scala 41:29]
  reg  way0_dirty_91; // @[data_cache.scala 41:29]
  reg  way0_dirty_92; // @[data_cache.scala 41:29]
  reg  way0_dirty_93; // @[data_cache.scala 41:29]
  reg  way0_dirty_94; // @[data_cache.scala 41:29]
  reg  way0_dirty_95; // @[data_cache.scala 41:29]
  reg  way0_dirty_96; // @[data_cache.scala 41:29]
  reg  way0_dirty_97; // @[data_cache.scala 41:29]
  reg  way0_dirty_98; // @[data_cache.scala 41:29]
  reg  way0_dirty_99; // @[data_cache.scala 41:29]
  reg  way0_dirty_100; // @[data_cache.scala 41:29]
  reg  way0_dirty_101; // @[data_cache.scala 41:29]
  reg  way0_dirty_102; // @[data_cache.scala 41:29]
  reg  way0_dirty_103; // @[data_cache.scala 41:29]
  reg  way0_dirty_104; // @[data_cache.scala 41:29]
  reg  way0_dirty_105; // @[data_cache.scala 41:29]
  reg  way0_dirty_106; // @[data_cache.scala 41:29]
  reg  way0_dirty_107; // @[data_cache.scala 41:29]
  reg  way0_dirty_108; // @[data_cache.scala 41:29]
  reg  way0_dirty_109; // @[data_cache.scala 41:29]
  reg  way0_dirty_110; // @[data_cache.scala 41:29]
  reg  way0_dirty_111; // @[data_cache.scala 41:29]
  reg  way0_dirty_112; // @[data_cache.scala 41:29]
  reg  way0_dirty_113; // @[data_cache.scala 41:29]
  reg  way0_dirty_114; // @[data_cache.scala 41:29]
  reg  way0_dirty_115; // @[data_cache.scala 41:29]
  reg  way0_dirty_116; // @[data_cache.scala 41:29]
  reg  way0_dirty_117; // @[data_cache.scala 41:29]
  reg  way0_dirty_118; // @[data_cache.scala 41:29]
  reg  way0_dirty_119; // @[data_cache.scala 41:29]
  reg  way0_dirty_120; // @[data_cache.scala 41:29]
  reg  way0_dirty_121; // @[data_cache.scala 41:29]
  reg  way0_dirty_122; // @[data_cache.scala 41:29]
  reg  way0_dirty_123; // @[data_cache.scala 41:29]
  reg  way0_dirty_124; // @[data_cache.scala 41:29]
  reg  way0_dirty_125; // @[data_cache.scala 41:29]
  reg  way0_dirty_126; // @[data_cache.scala 41:29]
  reg  way0_dirty_127; // @[data_cache.scala 41:29]
  reg  way1_dirty_0; // @[data_cache.scala 42:29]
  reg  way1_dirty_1; // @[data_cache.scala 42:29]
  reg  way1_dirty_2; // @[data_cache.scala 42:29]
  reg  way1_dirty_3; // @[data_cache.scala 42:29]
  reg  way1_dirty_4; // @[data_cache.scala 42:29]
  reg  way1_dirty_5; // @[data_cache.scala 42:29]
  reg  way1_dirty_6; // @[data_cache.scala 42:29]
  reg  way1_dirty_7; // @[data_cache.scala 42:29]
  reg  way1_dirty_8; // @[data_cache.scala 42:29]
  reg  way1_dirty_9; // @[data_cache.scala 42:29]
  reg  way1_dirty_10; // @[data_cache.scala 42:29]
  reg  way1_dirty_11; // @[data_cache.scala 42:29]
  reg  way1_dirty_12; // @[data_cache.scala 42:29]
  reg  way1_dirty_13; // @[data_cache.scala 42:29]
  reg  way1_dirty_14; // @[data_cache.scala 42:29]
  reg  way1_dirty_15; // @[data_cache.scala 42:29]
  reg  way1_dirty_16; // @[data_cache.scala 42:29]
  reg  way1_dirty_17; // @[data_cache.scala 42:29]
  reg  way1_dirty_18; // @[data_cache.scala 42:29]
  reg  way1_dirty_19; // @[data_cache.scala 42:29]
  reg  way1_dirty_20; // @[data_cache.scala 42:29]
  reg  way1_dirty_21; // @[data_cache.scala 42:29]
  reg  way1_dirty_22; // @[data_cache.scala 42:29]
  reg  way1_dirty_23; // @[data_cache.scala 42:29]
  reg  way1_dirty_24; // @[data_cache.scala 42:29]
  reg  way1_dirty_25; // @[data_cache.scala 42:29]
  reg  way1_dirty_26; // @[data_cache.scala 42:29]
  reg  way1_dirty_27; // @[data_cache.scala 42:29]
  reg  way1_dirty_28; // @[data_cache.scala 42:29]
  reg  way1_dirty_29; // @[data_cache.scala 42:29]
  reg  way1_dirty_30; // @[data_cache.scala 42:29]
  reg  way1_dirty_31; // @[data_cache.scala 42:29]
  reg  way1_dirty_32; // @[data_cache.scala 42:29]
  reg  way1_dirty_33; // @[data_cache.scala 42:29]
  reg  way1_dirty_34; // @[data_cache.scala 42:29]
  reg  way1_dirty_35; // @[data_cache.scala 42:29]
  reg  way1_dirty_36; // @[data_cache.scala 42:29]
  reg  way1_dirty_37; // @[data_cache.scala 42:29]
  reg  way1_dirty_38; // @[data_cache.scala 42:29]
  reg  way1_dirty_39; // @[data_cache.scala 42:29]
  reg  way1_dirty_40; // @[data_cache.scala 42:29]
  reg  way1_dirty_41; // @[data_cache.scala 42:29]
  reg  way1_dirty_42; // @[data_cache.scala 42:29]
  reg  way1_dirty_43; // @[data_cache.scala 42:29]
  reg  way1_dirty_44; // @[data_cache.scala 42:29]
  reg  way1_dirty_45; // @[data_cache.scala 42:29]
  reg  way1_dirty_46; // @[data_cache.scala 42:29]
  reg  way1_dirty_47; // @[data_cache.scala 42:29]
  reg  way1_dirty_48; // @[data_cache.scala 42:29]
  reg  way1_dirty_49; // @[data_cache.scala 42:29]
  reg  way1_dirty_50; // @[data_cache.scala 42:29]
  reg  way1_dirty_51; // @[data_cache.scala 42:29]
  reg  way1_dirty_52; // @[data_cache.scala 42:29]
  reg  way1_dirty_53; // @[data_cache.scala 42:29]
  reg  way1_dirty_54; // @[data_cache.scala 42:29]
  reg  way1_dirty_55; // @[data_cache.scala 42:29]
  reg  way1_dirty_56; // @[data_cache.scala 42:29]
  reg  way1_dirty_57; // @[data_cache.scala 42:29]
  reg  way1_dirty_58; // @[data_cache.scala 42:29]
  reg  way1_dirty_59; // @[data_cache.scala 42:29]
  reg  way1_dirty_60; // @[data_cache.scala 42:29]
  reg  way1_dirty_61; // @[data_cache.scala 42:29]
  reg  way1_dirty_62; // @[data_cache.scala 42:29]
  reg  way1_dirty_63; // @[data_cache.scala 42:29]
  reg  way1_dirty_64; // @[data_cache.scala 42:29]
  reg  way1_dirty_65; // @[data_cache.scala 42:29]
  reg  way1_dirty_66; // @[data_cache.scala 42:29]
  reg  way1_dirty_67; // @[data_cache.scala 42:29]
  reg  way1_dirty_68; // @[data_cache.scala 42:29]
  reg  way1_dirty_69; // @[data_cache.scala 42:29]
  reg  way1_dirty_70; // @[data_cache.scala 42:29]
  reg  way1_dirty_71; // @[data_cache.scala 42:29]
  reg  way1_dirty_72; // @[data_cache.scala 42:29]
  reg  way1_dirty_73; // @[data_cache.scala 42:29]
  reg  way1_dirty_74; // @[data_cache.scala 42:29]
  reg  way1_dirty_75; // @[data_cache.scala 42:29]
  reg  way1_dirty_76; // @[data_cache.scala 42:29]
  reg  way1_dirty_77; // @[data_cache.scala 42:29]
  reg  way1_dirty_78; // @[data_cache.scala 42:29]
  reg  way1_dirty_79; // @[data_cache.scala 42:29]
  reg  way1_dirty_80; // @[data_cache.scala 42:29]
  reg  way1_dirty_81; // @[data_cache.scala 42:29]
  reg  way1_dirty_82; // @[data_cache.scala 42:29]
  reg  way1_dirty_83; // @[data_cache.scala 42:29]
  reg  way1_dirty_84; // @[data_cache.scala 42:29]
  reg  way1_dirty_85; // @[data_cache.scala 42:29]
  reg  way1_dirty_86; // @[data_cache.scala 42:29]
  reg  way1_dirty_87; // @[data_cache.scala 42:29]
  reg  way1_dirty_88; // @[data_cache.scala 42:29]
  reg  way1_dirty_89; // @[data_cache.scala 42:29]
  reg  way1_dirty_90; // @[data_cache.scala 42:29]
  reg  way1_dirty_91; // @[data_cache.scala 42:29]
  reg  way1_dirty_92; // @[data_cache.scala 42:29]
  reg  way1_dirty_93; // @[data_cache.scala 42:29]
  reg  way1_dirty_94; // @[data_cache.scala 42:29]
  reg  way1_dirty_95; // @[data_cache.scala 42:29]
  reg  way1_dirty_96; // @[data_cache.scala 42:29]
  reg  way1_dirty_97; // @[data_cache.scala 42:29]
  reg  way1_dirty_98; // @[data_cache.scala 42:29]
  reg  way1_dirty_99; // @[data_cache.scala 42:29]
  reg  way1_dirty_100; // @[data_cache.scala 42:29]
  reg  way1_dirty_101; // @[data_cache.scala 42:29]
  reg  way1_dirty_102; // @[data_cache.scala 42:29]
  reg  way1_dirty_103; // @[data_cache.scala 42:29]
  reg  way1_dirty_104; // @[data_cache.scala 42:29]
  reg  way1_dirty_105; // @[data_cache.scala 42:29]
  reg  way1_dirty_106; // @[data_cache.scala 42:29]
  reg  way1_dirty_107; // @[data_cache.scala 42:29]
  reg  way1_dirty_108; // @[data_cache.scala 42:29]
  reg  way1_dirty_109; // @[data_cache.scala 42:29]
  reg  way1_dirty_110; // @[data_cache.scala 42:29]
  reg  way1_dirty_111; // @[data_cache.scala 42:29]
  reg  way1_dirty_112; // @[data_cache.scala 42:29]
  reg  way1_dirty_113; // @[data_cache.scala 42:29]
  reg  way1_dirty_114; // @[data_cache.scala 42:29]
  reg  way1_dirty_115; // @[data_cache.scala 42:29]
  reg  way1_dirty_116; // @[data_cache.scala 42:29]
  reg  way1_dirty_117; // @[data_cache.scala 42:29]
  reg  way1_dirty_118; // @[data_cache.scala 42:29]
  reg  way1_dirty_119; // @[data_cache.scala 42:29]
  reg  way1_dirty_120; // @[data_cache.scala 42:29]
  reg  way1_dirty_121; // @[data_cache.scala 42:29]
  reg  way1_dirty_122; // @[data_cache.scala 42:29]
  reg  way1_dirty_123; // @[data_cache.scala 42:29]
  reg  way1_dirty_124; // @[data_cache.scala 42:29]
  reg  way1_dirty_125; // @[data_cache.scala 42:29]
  reg  way1_dirty_126; // @[data_cache.scala 42:29]
  reg  way1_dirty_127; // @[data_cache.scala 42:29]
  reg [31:0] stage1_sram_addr_reg; // @[data_cache.scala 46:39]
  reg  stage1_sram_cache_reg; // @[data_cache.scala 47:40]
  reg [31:0] stage1_sram_wdata_reg; // @[data_cache.scala 48:40]
  reg [1:0] stage1_sram_size_reg; // @[data_cache.scala 49:39]
  reg  stage1_sram_wr_reg; // @[data_cache.scala 50:37]
  reg  stage1_sram_req_reg; // @[data_cache.scala 51:38]
  reg  stage1_sram_hit0_reg; // @[data_cache.scala 53:40]
  reg  stage1_sram_hit1_reg; // @[data_cache.scala 54:40]
  reg  stage1_sram_valid0_reg; // @[data_cache.scala 55:42]
  reg  stage1_sram_valid1_reg; // @[data_cache.scala 56:42]
  reg [3:0] stage1_wstrb_reg; // @[data_cache.scala 57:35]
  reg [31:0] stage1_sram_phy_addr_reg; // @[data_cache.scala 59:43]
  reg [2:0] stage1_exception; // @[data_cache.scala 60:37]
  wire  _hit_T = stage1_sram_hit0_reg & stage1_sram_valid0_reg; // @[data_cache.scala 185:37]
  wire  _hit_T_1 = stage1_sram_hit1_reg & stage1_sram_valid1_reg; // @[data_cache.scala 186:31]
  wire  hit = stage1_sram_hit0_reg & stage1_sram_valid0_reg | _hit_T_1; // @[data_cache.scala 185:64]
  wire [4:0] _state_ready_lookup_should_be_T_2 = stage1_sram_cache_reg ? 5'h19 : 5'h0; // @[data_cache.scala 194:82]
  wire [4:0] _state_ready_lookup_should_be_T_3 = stage1_sram_req_reg ? _state_ready_lookup_should_be_T_2 : 5'h19; // @[data_cache.scala 194:51]
  wire [4:0] _state_ready_lookup_should_be_T_5 = stage1_sram_req_reg ? 5'h0 : 5'h19; // @[data_cache.scala 195:16]
  wire [4:0] state_ready_lookup_should_be = hit ? _state_ready_lookup_should_be_T_3 : _state_ready_lookup_should_be_T_5; // @[data_cache.scala 194:43]
  wire [4:0] _access_work_state_for_stall_T_1 = io_port_rvalid ? 5'h18 : work_state; // @[data_cache.scala 221:39]
  wire [4:0] _access_work_state_for_stall_T_3 = 5'h2 == work_state ? _access_work_state_for_stall_T_1 : work_state; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_for_stall_T_5 = 5'h18 == work_state ? state_ready_lookup_should_be :
    _access_work_state_for_stall_T_3; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_for_stall_T_7 = 5'h5 == work_state ? 5'h18 : _access_work_state_for_stall_T_5; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_for_stall_T_9 = 5'h19 == work_state ? state_ready_lookup_should_be :
    _access_work_state_for_stall_T_7; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_for_stall_T_11 = 5'he == work_state ? 5'h18 : _access_work_state_for_stall_T_9; // @[Mux.scala 81:58]
  wire [4:0] access_work_state_for_stall = 5'h10 == work_state ? 5'h18 : _access_work_state_for_stall_T_11; // @[Mux.scala 81:58]
  wire  _stage2_stall_T_2 = stage1_exception != 3'h0; // @[data_cache.scala 232:86]
  wire  stage2_stall = access_work_state_for_stall[4:3] == 2'h3 | stage1_exception != 3'h0; // @[data_cache.scala 232:66]
  reg  stage2_sram_write_reg; // @[data_cache.scala 123:40]
  reg  stage1_stall_reg; // @[data_cache.scala 130:35]
  reg  write_access_complete_reg; // @[data_cache.scala 133:44]
  wire  _stage1_sram_req_reg_T_1 = stage2_stall ? 1'h0 : stage1_sram_req_reg; // @[data_cache.scala 142:65]
  wire [4:0] _state_lookup_for_less_delay_T_1 = 5'h18 == work_state ? state_ready_lookup_should_be : work_state; // @[Mux.scala 81:58]
  wire [4:0] state_lookup_for_less_delay = 5'h19 == work_state ? state_ready_lookup_should_be :
    _state_lookup_for_less_delay_T_1; // @[Mux.scala 81:58]
  wire  _way0_dirty_T = state_lookup_for_less_delay == 5'h19; // @[data_cache.scala 151:79]
  wire  _way0_dirty_T_2 = state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg; // @[data_cache.scala 151:96]
  wire  _way0_dirty_T_4 = state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
    stage1_sram_valid0_reg; // @[data_cache.scala 151:149]
  wire  _way0_dirty_T_5 = work_state == 5'he; // @[data_cache.scala 152:24]
  wire  _GEN_2 = 7'h1 == stage1_sram_addr_reg[11:5] ? lru_1 : lru_0; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_3 = 7'h2 == stage1_sram_addr_reg[11:5] ? lru_2 : _GEN_2; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_4 = 7'h3 == stage1_sram_addr_reg[11:5] ? lru_3 : _GEN_3; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_5 = 7'h4 == stage1_sram_addr_reg[11:5] ? lru_4 : _GEN_4; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_6 = 7'h5 == stage1_sram_addr_reg[11:5] ? lru_5 : _GEN_5; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_7 = 7'h6 == stage1_sram_addr_reg[11:5] ? lru_6 : _GEN_6; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_8 = 7'h7 == stage1_sram_addr_reg[11:5] ? lru_7 : _GEN_7; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_9 = 7'h8 == stage1_sram_addr_reg[11:5] ? lru_8 : _GEN_8; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_10 = 7'h9 == stage1_sram_addr_reg[11:5] ? lru_9 : _GEN_9; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_11 = 7'ha == stage1_sram_addr_reg[11:5] ? lru_10 : _GEN_10; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_12 = 7'hb == stage1_sram_addr_reg[11:5] ? lru_11 : _GEN_11; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_13 = 7'hc == stage1_sram_addr_reg[11:5] ? lru_12 : _GEN_12; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_14 = 7'hd == stage1_sram_addr_reg[11:5] ? lru_13 : _GEN_13; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_15 = 7'he == stage1_sram_addr_reg[11:5] ? lru_14 : _GEN_14; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_16 = 7'hf == stage1_sram_addr_reg[11:5] ? lru_15 : _GEN_15; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_17 = 7'h10 == stage1_sram_addr_reg[11:5] ? lru_16 : _GEN_16; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_18 = 7'h11 == stage1_sram_addr_reg[11:5] ? lru_17 : _GEN_17; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_19 = 7'h12 == stage1_sram_addr_reg[11:5] ? lru_18 : _GEN_18; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_20 = 7'h13 == stage1_sram_addr_reg[11:5] ? lru_19 : _GEN_19; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_21 = 7'h14 == stage1_sram_addr_reg[11:5] ? lru_20 : _GEN_20; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_22 = 7'h15 == stage1_sram_addr_reg[11:5] ? lru_21 : _GEN_21; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_23 = 7'h16 == stage1_sram_addr_reg[11:5] ? lru_22 : _GEN_22; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_24 = 7'h17 == stage1_sram_addr_reg[11:5] ? lru_23 : _GEN_23; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_25 = 7'h18 == stage1_sram_addr_reg[11:5] ? lru_24 : _GEN_24; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_26 = 7'h19 == stage1_sram_addr_reg[11:5] ? lru_25 : _GEN_25; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_27 = 7'h1a == stage1_sram_addr_reg[11:5] ? lru_26 : _GEN_26; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_28 = 7'h1b == stage1_sram_addr_reg[11:5] ? lru_27 : _GEN_27; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_29 = 7'h1c == stage1_sram_addr_reg[11:5] ? lru_28 : _GEN_28; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_30 = 7'h1d == stage1_sram_addr_reg[11:5] ? lru_29 : _GEN_29; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_31 = 7'h1e == stage1_sram_addr_reg[11:5] ? lru_30 : _GEN_30; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_32 = 7'h1f == stage1_sram_addr_reg[11:5] ? lru_31 : _GEN_31; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_33 = 7'h20 == stage1_sram_addr_reg[11:5] ? lru_32 : _GEN_32; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_34 = 7'h21 == stage1_sram_addr_reg[11:5] ? lru_33 : _GEN_33; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_35 = 7'h22 == stage1_sram_addr_reg[11:5] ? lru_34 : _GEN_34; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_36 = 7'h23 == stage1_sram_addr_reg[11:5] ? lru_35 : _GEN_35; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_37 = 7'h24 == stage1_sram_addr_reg[11:5] ? lru_36 : _GEN_36; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_38 = 7'h25 == stage1_sram_addr_reg[11:5] ? lru_37 : _GEN_37; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_39 = 7'h26 == stage1_sram_addr_reg[11:5] ? lru_38 : _GEN_38; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_40 = 7'h27 == stage1_sram_addr_reg[11:5] ? lru_39 : _GEN_39; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_41 = 7'h28 == stage1_sram_addr_reg[11:5] ? lru_40 : _GEN_40; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_42 = 7'h29 == stage1_sram_addr_reg[11:5] ? lru_41 : _GEN_41; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_43 = 7'h2a == stage1_sram_addr_reg[11:5] ? lru_42 : _GEN_42; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_44 = 7'h2b == stage1_sram_addr_reg[11:5] ? lru_43 : _GEN_43; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_45 = 7'h2c == stage1_sram_addr_reg[11:5] ? lru_44 : _GEN_44; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_46 = 7'h2d == stage1_sram_addr_reg[11:5] ? lru_45 : _GEN_45; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_47 = 7'h2e == stage1_sram_addr_reg[11:5] ? lru_46 : _GEN_46; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_48 = 7'h2f == stage1_sram_addr_reg[11:5] ? lru_47 : _GEN_47; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_49 = 7'h30 == stage1_sram_addr_reg[11:5] ? lru_48 : _GEN_48; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_50 = 7'h31 == stage1_sram_addr_reg[11:5] ? lru_49 : _GEN_49; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_51 = 7'h32 == stage1_sram_addr_reg[11:5] ? lru_50 : _GEN_50; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_52 = 7'h33 == stage1_sram_addr_reg[11:5] ? lru_51 : _GEN_51; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_53 = 7'h34 == stage1_sram_addr_reg[11:5] ? lru_52 : _GEN_52; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_54 = 7'h35 == stage1_sram_addr_reg[11:5] ? lru_53 : _GEN_53; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_55 = 7'h36 == stage1_sram_addr_reg[11:5] ? lru_54 : _GEN_54; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_56 = 7'h37 == stage1_sram_addr_reg[11:5] ? lru_55 : _GEN_55; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_57 = 7'h38 == stage1_sram_addr_reg[11:5] ? lru_56 : _GEN_56; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_58 = 7'h39 == stage1_sram_addr_reg[11:5] ? lru_57 : _GEN_57; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_59 = 7'h3a == stage1_sram_addr_reg[11:5] ? lru_58 : _GEN_58; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_60 = 7'h3b == stage1_sram_addr_reg[11:5] ? lru_59 : _GEN_59; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_61 = 7'h3c == stage1_sram_addr_reg[11:5] ? lru_60 : _GEN_60; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_62 = 7'h3d == stage1_sram_addr_reg[11:5] ? lru_61 : _GEN_61; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_63 = 7'h3e == stage1_sram_addr_reg[11:5] ? lru_62 : _GEN_62; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_64 = 7'h3f == stage1_sram_addr_reg[11:5] ? lru_63 : _GEN_63; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_65 = 7'h40 == stage1_sram_addr_reg[11:5] ? lru_64 : _GEN_64; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_66 = 7'h41 == stage1_sram_addr_reg[11:5] ? lru_65 : _GEN_65; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_67 = 7'h42 == stage1_sram_addr_reg[11:5] ? lru_66 : _GEN_66; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_68 = 7'h43 == stage1_sram_addr_reg[11:5] ? lru_67 : _GEN_67; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_69 = 7'h44 == stage1_sram_addr_reg[11:5] ? lru_68 : _GEN_68; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_70 = 7'h45 == stage1_sram_addr_reg[11:5] ? lru_69 : _GEN_69; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_71 = 7'h46 == stage1_sram_addr_reg[11:5] ? lru_70 : _GEN_70; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_72 = 7'h47 == stage1_sram_addr_reg[11:5] ? lru_71 : _GEN_71; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_73 = 7'h48 == stage1_sram_addr_reg[11:5] ? lru_72 : _GEN_72; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_74 = 7'h49 == stage1_sram_addr_reg[11:5] ? lru_73 : _GEN_73; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_75 = 7'h4a == stage1_sram_addr_reg[11:5] ? lru_74 : _GEN_74; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_76 = 7'h4b == stage1_sram_addr_reg[11:5] ? lru_75 : _GEN_75; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_77 = 7'h4c == stage1_sram_addr_reg[11:5] ? lru_76 : _GEN_76; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_78 = 7'h4d == stage1_sram_addr_reg[11:5] ? lru_77 : _GEN_77; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_79 = 7'h4e == stage1_sram_addr_reg[11:5] ? lru_78 : _GEN_78; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_80 = 7'h4f == stage1_sram_addr_reg[11:5] ? lru_79 : _GEN_79; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_81 = 7'h50 == stage1_sram_addr_reg[11:5] ? lru_80 : _GEN_80; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_82 = 7'h51 == stage1_sram_addr_reg[11:5] ? lru_81 : _GEN_81; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_83 = 7'h52 == stage1_sram_addr_reg[11:5] ? lru_82 : _GEN_82; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_84 = 7'h53 == stage1_sram_addr_reg[11:5] ? lru_83 : _GEN_83; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_85 = 7'h54 == stage1_sram_addr_reg[11:5] ? lru_84 : _GEN_84; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_86 = 7'h55 == stage1_sram_addr_reg[11:5] ? lru_85 : _GEN_85; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_87 = 7'h56 == stage1_sram_addr_reg[11:5] ? lru_86 : _GEN_86; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_88 = 7'h57 == stage1_sram_addr_reg[11:5] ? lru_87 : _GEN_87; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_89 = 7'h58 == stage1_sram_addr_reg[11:5] ? lru_88 : _GEN_88; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_90 = 7'h59 == stage1_sram_addr_reg[11:5] ? lru_89 : _GEN_89; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_91 = 7'h5a == stage1_sram_addr_reg[11:5] ? lru_90 : _GEN_90; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_92 = 7'h5b == stage1_sram_addr_reg[11:5] ? lru_91 : _GEN_91; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_93 = 7'h5c == stage1_sram_addr_reg[11:5] ? lru_92 : _GEN_92; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_94 = 7'h5d == stage1_sram_addr_reg[11:5] ? lru_93 : _GEN_93; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_95 = 7'h5e == stage1_sram_addr_reg[11:5] ? lru_94 : _GEN_94; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_96 = 7'h5f == stage1_sram_addr_reg[11:5] ? lru_95 : _GEN_95; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_97 = 7'h60 == stage1_sram_addr_reg[11:5] ? lru_96 : _GEN_96; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_98 = 7'h61 == stage1_sram_addr_reg[11:5] ? lru_97 : _GEN_97; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_99 = 7'h62 == stage1_sram_addr_reg[11:5] ? lru_98 : _GEN_98; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_100 = 7'h63 == stage1_sram_addr_reg[11:5] ? lru_99 : _GEN_99; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_101 = 7'h64 == stage1_sram_addr_reg[11:5] ? lru_100 : _GEN_100; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_102 = 7'h65 == stage1_sram_addr_reg[11:5] ? lru_101 : _GEN_101; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_103 = 7'h66 == stage1_sram_addr_reg[11:5] ? lru_102 : _GEN_102; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_104 = 7'h67 == stage1_sram_addr_reg[11:5] ? lru_103 : _GEN_103; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_105 = 7'h68 == stage1_sram_addr_reg[11:5] ? lru_104 : _GEN_104; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_106 = 7'h69 == stage1_sram_addr_reg[11:5] ? lru_105 : _GEN_105; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_107 = 7'h6a == stage1_sram_addr_reg[11:5] ? lru_106 : _GEN_106; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_108 = 7'h6b == stage1_sram_addr_reg[11:5] ? lru_107 : _GEN_107; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_109 = 7'h6c == stage1_sram_addr_reg[11:5] ? lru_108 : _GEN_108; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_110 = 7'h6d == stage1_sram_addr_reg[11:5] ? lru_109 : _GEN_109; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_111 = 7'h6e == stage1_sram_addr_reg[11:5] ? lru_110 : _GEN_110; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_112 = 7'h6f == stage1_sram_addr_reg[11:5] ? lru_111 : _GEN_111; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_113 = 7'h70 == stage1_sram_addr_reg[11:5] ? lru_112 : _GEN_112; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_114 = 7'h71 == stage1_sram_addr_reg[11:5] ? lru_113 : _GEN_113; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_115 = 7'h72 == stage1_sram_addr_reg[11:5] ? lru_114 : _GEN_114; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_116 = 7'h73 == stage1_sram_addr_reg[11:5] ? lru_115 : _GEN_115; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_117 = 7'h74 == stage1_sram_addr_reg[11:5] ? lru_116 : _GEN_116; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_118 = 7'h75 == stage1_sram_addr_reg[11:5] ? lru_117 : _GEN_117; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_119 = 7'h76 == stage1_sram_addr_reg[11:5] ? lru_118 : _GEN_118; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_120 = 7'h77 == stage1_sram_addr_reg[11:5] ? lru_119 : _GEN_119; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_121 = 7'h78 == stage1_sram_addr_reg[11:5] ? lru_120 : _GEN_120; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_122 = 7'h79 == stage1_sram_addr_reg[11:5] ? lru_121 : _GEN_121; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_123 = 7'h7a == stage1_sram_addr_reg[11:5] ? lru_122 : _GEN_122; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_124 = 7'h7b == stage1_sram_addr_reg[11:5] ? lru_123 : _GEN_123; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_125 = 7'h7c == stage1_sram_addr_reg[11:5] ? lru_124 : _GEN_124; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_126 = 7'h7d == stage1_sram_addr_reg[11:5] ? lru_125 : _GEN_125; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_127 = 7'h7e == stage1_sram_addr_reg[11:5] ? lru_126 : _GEN_126; // @[data_cache.scala 152:{86,86}]
  wire  _GEN_128 = 7'h7f == stage1_sram_addr_reg[11:5] ? lru_127 : _GEN_127; // @[data_cache.scala 152:{86,86}]
  wire  _way0_dirty_T_7 = ~_GEN_128; // @[data_cache.scala 152:86]
  wire  _way0_dirty_T_9 = work_state == 5'h10; // @[data_cache.scala 153:24]
  wire  _way0_dirty_T_12 = work_state == 5'h10 & _way0_dirty_T_7; // @[data_cache.scala 153:52]
  wire  _GEN_258 = 7'h1 == stage1_sram_addr_reg[11:5] ? way0_dirty_1 : way0_dirty_0; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_259 = 7'h2 == stage1_sram_addr_reg[11:5] ? way0_dirty_2 : _GEN_258; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_260 = 7'h3 == stage1_sram_addr_reg[11:5] ? way0_dirty_3 : _GEN_259; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_261 = 7'h4 == stage1_sram_addr_reg[11:5] ? way0_dirty_4 : _GEN_260; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_262 = 7'h5 == stage1_sram_addr_reg[11:5] ? way0_dirty_5 : _GEN_261; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_263 = 7'h6 == stage1_sram_addr_reg[11:5] ? way0_dirty_6 : _GEN_262; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_264 = 7'h7 == stage1_sram_addr_reg[11:5] ? way0_dirty_7 : _GEN_263; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_265 = 7'h8 == stage1_sram_addr_reg[11:5] ? way0_dirty_8 : _GEN_264; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_266 = 7'h9 == stage1_sram_addr_reg[11:5] ? way0_dirty_9 : _GEN_265; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_267 = 7'ha == stage1_sram_addr_reg[11:5] ? way0_dirty_10 : _GEN_266; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_268 = 7'hb == stage1_sram_addr_reg[11:5] ? way0_dirty_11 : _GEN_267; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_269 = 7'hc == stage1_sram_addr_reg[11:5] ? way0_dirty_12 : _GEN_268; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_270 = 7'hd == stage1_sram_addr_reg[11:5] ? way0_dirty_13 : _GEN_269; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_271 = 7'he == stage1_sram_addr_reg[11:5] ? way0_dirty_14 : _GEN_270; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_272 = 7'hf == stage1_sram_addr_reg[11:5] ? way0_dirty_15 : _GEN_271; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_273 = 7'h10 == stage1_sram_addr_reg[11:5] ? way0_dirty_16 : _GEN_272; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_274 = 7'h11 == stage1_sram_addr_reg[11:5] ? way0_dirty_17 : _GEN_273; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_275 = 7'h12 == stage1_sram_addr_reg[11:5] ? way0_dirty_18 : _GEN_274; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_276 = 7'h13 == stage1_sram_addr_reg[11:5] ? way0_dirty_19 : _GEN_275; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_277 = 7'h14 == stage1_sram_addr_reg[11:5] ? way0_dirty_20 : _GEN_276; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_278 = 7'h15 == stage1_sram_addr_reg[11:5] ? way0_dirty_21 : _GEN_277; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_279 = 7'h16 == stage1_sram_addr_reg[11:5] ? way0_dirty_22 : _GEN_278; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_280 = 7'h17 == stage1_sram_addr_reg[11:5] ? way0_dirty_23 : _GEN_279; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_281 = 7'h18 == stage1_sram_addr_reg[11:5] ? way0_dirty_24 : _GEN_280; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_282 = 7'h19 == stage1_sram_addr_reg[11:5] ? way0_dirty_25 : _GEN_281; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_283 = 7'h1a == stage1_sram_addr_reg[11:5] ? way0_dirty_26 : _GEN_282; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_284 = 7'h1b == stage1_sram_addr_reg[11:5] ? way0_dirty_27 : _GEN_283; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_285 = 7'h1c == stage1_sram_addr_reg[11:5] ? way0_dirty_28 : _GEN_284; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_286 = 7'h1d == stage1_sram_addr_reg[11:5] ? way0_dirty_29 : _GEN_285; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_287 = 7'h1e == stage1_sram_addr_reg[11:5] ? way0_dirty_30 : _GEN_286; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_288 = 7'h1f == stage1_sram_addr_reg[11:5] ? way0_dirty_31 : _GEN_287; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_289 = 7'h20 == stage1_sram_addr_reg[11:5] ? way0_dirty_32 : _GEN_288; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_290 = 7'h21 == stage1_sram_addr_reg[11:5] ? way0_dirty_33 : _GEN_289; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_291 = 7'h22 == stage1_sram_addr_reg[11:5] ? way0_dirty_34 : _GEN_290; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_292 = 7'h23 == stage1_sram_addr_reg[11:5] ? way0_dirty_35 : _GEN_291; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_293 = 7'h24 == stage1_sram_addr_reg[11:5] ? way0_dirty_36 : _GEN_292; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_294 = 7'h25 == stage1_sram_addr_reg[11:5] ? way0_dirty_37 : _GEN_293; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_295 = 7'h26 == stage1_sram_addr_reg[11:5] ? way0_dirty_38 : _GEN_294; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_296 = 7'h27 == stage1_sram_addr_reg[11:5] ? way0_dirty_39 : _GEN_295; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_297 = 7'h28 == stage1_sram_addr_reg[11:5] ? way0_dirty_40 : _GEN_296; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_298 = 7'h29 == stage1_sram_addr_reg[11:5] ? way0_dirty_41 : _GEN_297; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_299 = 7'h2a == stage1_sram_addr_reg[11:5] ? way0_dirty_42 : _GEN_298; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_300 = 7'h2b == stage1_sram_addr_reg[11:5] ? way0_dirty_43 : _GEN_299; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_301 = 7'h2c == stage1_sram_addr_reg[11:5] ? way0_dirty_44 : _GEN_300; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_302 = 7'h2d == stage1_sram_addr_reg[11:5] ? way0_dirty_45 : _GEN_301; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_303 = 7'h2e == stage1_sram_addr_reg[11:5] ? way0_dirty_46 : _GEN_302; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_304 = 7'h2f == stage1_sram_addr_reg[11:5] ? way0_dirty_47 : _GEN_303; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_305 = 7'h30 == stage1_sram_addr_reg[11:5] ? way0_dirty_48 : _GEN_304; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_306 = 7'h31 == stage1_sram_addr_reg[11:5] ? way0_dirty_49 : _GEN_305; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_307 = 7'h32 == stage1_sram_addr_reg[11:5] ? way0_dirty_50 : _GEN_306; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_308 = 7'h33 == stage1_sram_addr_reg[11:5] ? way0_dirty_51 : _GEN_307; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_309 = 7'h34 == stage1_sram_addr_reg[11:5] ? way0_dirty_52 : _GEN_308; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_310 = 7'h35 == stage1_sram_addr_reg[11:5] ? way0_dirty_53 : _GEN_309; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_311 = 7'h36 == stage1_sram_addr_reg[11:5] ? way0_dirty_54 : _GEN_310; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_312 = 7'h37 == stage1_sram_addr_reg[11:5] ? way0_dirty_55 : _GEN_311; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_313 = 7'h38 == stage1_sram_addr_reg[11:5] ? way0_dirty_56 : _GEN_312; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_314 = 7'h39 == stage1_sram_addr_reg[11:5] ? way0_dirty_57 : _GEN_313; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_315 = 7'h3a == stage1_sram_addr_reg[11:5] ? way0_dirty_58 : _GEN_314; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_316 = 7'h3b == stage1_sram_addr_reg[11:5] ? way0_dirty_59 : _GEN_315; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_317 = 7'h3c == stage1_sram_addr_reg[11:5] ? way0_dirty_60 : _GEN_316; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_318 = 7'h3d == stage1_sram_addr_reg[11:5] ? way0_dirty_61 : _GEN_317; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_319 = 7'h3e == stage1_sram_addr_reg[11:5] ? way0_dirty_62 : _GEN_318; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_320 = 7'h3f == stage1_sram_addr_reg[11:5] ? way0_dirty_63 : _GEN_319; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_321 = 7'h40 == stage1_sram_addr_reg[11:5] ? way0_dirty_64 : _GEN_320; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_322 = 7'h41 == stage1_sram_addr_reg[11:5] ? way0_dirty_65 : _GEN_321; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_323 = 7'h42 == stage1_sram_addr_reg[11:5] ? way0_dirty_66 : _GEN_322; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_324 = 7'h43 == stage1_sram_addr_reg[11:5] ? way0_dirty_67 : _GEN_323; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_325 = 7'h44 == stage1_sram_addr_reg[11:5] ? way0_dirty_68 : _GEN_324; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_326 = 7'h45 == stage1_sram_addr_reg[11:5] ? way0_dirty_69 : _GEN_325; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_327 = 7'h46 == stage1_sram_addr_reg[11:5] ? way0_dirty_70 : _GEN_326; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_328 = 7'h47 == stage1_sram_addr_reg[11:5] ? way0_dirty_71 : _GEN_327; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_329 = 7'h48 == stage1_sram_addr_reg[11:5] ? way0_dirty_72 : _GEN_328; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_330 = 7'h49 == stage1_sram_addr_reg[11:5] ? way0_dirty_73 : _GEN_329; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_331 = 7'h4a == stage1_sram_addr_reg[11:5] ? way0_dirty_74 : _GEN_330; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_332 = 7'h4b == stage1_sram_addr_reg[11:5] ? way0_dirty_75 : _GEN_331; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_333 = 7'h4c == stage1_sram_addr_reg[11:5] ? way0_dirty_76 : _GEN_332; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_334 = 7'h4d == stage1_sram_addr_reg[11:5] ? way0_dirty_77 : _GEN_333; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_335 = 7'h4e == stage1_sram_addr_reg[11:5] ? way0_dirty_78 : _GEN_334; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_336 = 7'h4f == stage1_sram_addr_reg[11:5] ? way0_dirty_79 : _GEN_335; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_337 = 7'h50 == stage1_sram_addr_reg[11:5] ? way0_dirty_80 : _GEN_336; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_338 = 7'h51 == stage1_sram_addr_reg[11:5] ? way0_dirty_81 : _GEN_337; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_339 = 7'h52 == stage1_sram_addr_reg[11:5] ? way0_dirty_82 : _GEN_338; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_340 = 7'h53 == stage1_sram_addr_reg[11:5] ? way0_dirty_83 : _GEN_339; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_341 = 7'h54 == stage1_sram_addr_reg[11:5] ? way0_dirty_84 : _GEN_340; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_342 = 7'h55 == stage1_sram_addr_reg[11:5] ? way0_dirty_85 : _GEN_341; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_343 = 7'h56 == stage1_sram_addr_reg[11:5] ? way0_dirty_86 : _GEN_342; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_344 = 7'h57 == stage1_sram_addr_reg[11:5] ? way0_dirty_87 : _GEN_343; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_345 = 7'h58 == stage1_sram_addr_reg[11:5] ? way0_dirty_88 : _GEN_344; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_346 = 7'h59 == stage1_sram_addr_reg[11:5] ? way0_dirty_89 : _GEN_345; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_347 = 7'h5a == stage1_sram_addr_reg[11:5] ? way0_dirty_90 : _GEN_346; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_348 = 7'h5b == stage1_sram_addr_reg[11:5] ? way0_dirty_91 : _GEN_347; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_349 = 7'h5c == stage1_sram_addr_reg[11:5] ? way0_dirty_92 : _GEN_348; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_350 = 7'h5d == stage1_sram_addr_reg[11:5] ? way0_dirty_93 : _GEN_349; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_351 = 7'h5e == stage1_sram_addr_reg[11:5] ? way0_dirty_94 : _GEN_350; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_352 = 7'h5f == stage1_sram_addr_reg[11:5] ? way0_dirty_95 : _GEN_351; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_353 = 7'h60 == stage1_sram_addr_reg[11:5] ? way0_dirty_96 : _GEN_352; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_354 = 7'h61 == stage1_sram_addr_reg[11:5] ? way0_dirty_97 : _GEN_353; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_355 = 7'h62 == stage1_sram_addr_reg[11:5] ? way0_dirty_98 : _GEN_354; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_356 = 7'h63 == stage1_sram_addr_reg[11:5] ? way0_dirty_99 : _GEN_355; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_357 = 7'h64 == stage1_sram_addr_reg[11:5] ? way0_dirty_100 : _GEN_356; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_358 = 7'h65 == stage1_sram_addr_reg[11:5] ? way0_dirty_101 : _GEN_357; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_359 = 7'h66 == stage1_sram_addr_reg[11:5] ? way0_dirty_102 : _GEN_358; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_360 = 7'h67 == stage1_sram_addr_reg[11:5] ? way0_dirty_103 : _GEN_359; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_361 = 7'h68 == stage1_sram_addr_reg[11:5] ? way0_dirty_104 : _GEN_360; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_362 = 7'h69 == stage1_sram_addr_reg[11:5] ? way0_dirty_105 : _GEN_361; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_363 = 7'h6a == stage1_sram_addr_reg[11:5] ? way0_dirty_106 : _GEN_362; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_364 = 7'h6b == stage1_sram_addr_reg[11:5] ? way0_dirty_107 : _GEN_363; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_365 = 7'h6c == stage1_sram_addr_reg[11:5] ? way0_dirty_108 : _GEN_364; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_366 = 7'h6d == stage1_sram_addr_reg[11:5] ? way0_dirty_109 : _GEN_365; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_367 = 7'h6e == stage1_sram_addr_reg[11:5] ? way0_dirty_110 : _GEN_366; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_368 = 7'h6f == stage1_sram_addr_reg[11:5] ? way0_dirty_111 : _GEN_367; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_369 = 7'h70 == stage1_sram_addr_reg[11:5] ? way0_dirty_112 : _GEN_368; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_370 = 7'h71 == stage1_sram_addr_reg[11:5] ? way0_dirty_113 : _GEN_369; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_371 = 7'h72 == stage1_sram_addr_reg[11:5] ? way0_dirty_114 : _GEN_370; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_372 = 7'h73 == stage1_sram_addr_reg[11:5] ? way0_dirty_115 : _GEN_371; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_373 = 7'h74 == stage1_sram_addr_reg[11:5] ? way0_dirty_116 : _GEN_372; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_374 = 7'h75 == stage1_sram_addr_reg[11:5] ? way0_dirty_117 : _GEN_373; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_375 = 7'h76 == stage1_sram_addr_reg[11:5] ? way0_dirty_118 : _GEN_374; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_376 = 7'h77 == stage1_sram_addr_reg[11:5] ? way0_dirty_119 : _GEN_375; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_377 = 7'h78 == stage1_sram_addr_reg[11:5] ? way0_dirty_120 : _GEN_376; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_378 = 7'h79 == stage1_sram_addr_reg[11:5] ? way0_dirty_121 : _GEN_377; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_379 = 7'h7a == stage1_sram_addr_reg[11:5] ? way0_dirty_122 : _GEN_378; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_380 = 7'h7b == stage1_sram_addr_reg[11:5] ? way0_dirty_123 : _GEN_379; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_381 = 7'h7c == stage1_sram_addr_reg[11:5] ? way0_dirty_124 : _GEN_380; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_382 = 7'h7d == stage1_sram_addr_reg[11:5] ? way0_dirty_125 : _GEN_381; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_383 = 7'h7e == stage1_sram_addr_reg[11:5] ? way0_dirty_126 : _GEN_382; // @[data_cache.scala 153:{12,12}]
  wire  _GEN_384 = 7'h7f == stage1_sram_addr_reg[11:5] ? way0_dirty_127 : _GEN_383; // @[data_cache.scala 153:{12,12}]
  wire  _way0_dirty_T_14 = work_state == 5'h10 & _way0_dirty_T_7 | _GEN_384; // @[data_cache.scala 153:12]
  wire  _way0_dirty_T_15 = work_state == 5'he & ~_GEN_128 ? 1'h0 : _way0_dirty_T_14; // @[data_cache.scala 152:12]
  wire  _way1_dirty_T_4 = _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg; // @[data_cache.scala 155:149]
  wire  _way1_dirty_T_12 = _way0_dirty_T_9 & _GEN_128; // @[data_cache.scala 157:52]
  wire  _GEN_770 = 7'h1 == stage1_sram_addr_reg[11:5] ? way1_dirty_1 : way1_dirty_0; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_771 = 7'h2 == stage1_sram_addr_reg[11:5] ? way1_dirty_2 : _GEN_770; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_772 = 7'h3 == stage1_sram_addr_reg[11:5] ? way1_dirty_3 : _GEN_771; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_773 = 7'h4 == stage1_sram_addr_reg[11:5] ? way1_dirty_4 : _GEN_772; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_774 = 7'h5 == stage1_sram_addr_reg[11:5] ? way1_dirty_5 : _GEN_773; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_775 = 7'h6 == stage1_sram_addr_reg[11:5] ? way1_dirty_6 : _GEN_774; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_776 = 7'h7 == stage1_sram_addr_reg[11:5] ? way1_dirty_7 : _GEN_775; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_777 = 7'h8 == stage1_sram_addr_reg[11:5] ? way1_dirty_8 : _GEN_776; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_778 = 7'h9 == stage1_sram_addr_reg[11:5] ? way1_dirty_9 : _GEN_777; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_779 = 7'ha == stage1_sram_addr_reg[11:5] ? way1_dirty_10 : _GEN_778; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_780 = 7'hb == stage1_sram_addr_reg[11:5] ? way1_dirty_11 : _GEN_779; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_781 = 7'hc == stage1_sram_addr_reg[11:5] ? way1_dirty_12 : _GEN_780; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_782 = 7'hd == stage1_sram_addr_reg[11:5] ? way1_dirty_13 : _GEN_781; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_783 = 7'he == stage1_sram_addr_reg[11:5] ? way1_dirty_14 : _GEN_782; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_784 = 7'hf == stage1_sram_addr_reg[11:5] ? way1_dirty_15 : _GEN_783; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_785 = 7'h10 == stage1_sram_addr_reg[11:5] ? way1_dirty_16 : _GEN_784; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_786 = 7'h11 == stage1_sram_addr_reg[11:5] ? way1_dirty_17 : _GEN_785; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_787 = 7'h12 == stage1_sram_addr_reg[11:5] ? way1_dirty_18 : _GEN_786; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_788 = 7'h13 == stage1_sram_addr_reg[11:5] ? way1_dirty_19 : _GEN_787; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_789 = 7'h14 == stage1_sram_addr_reg[11:5] ? way1_dirty_20 : _GEN_788; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_790 = 7'h15 == stage1_sram_addr_reg[11:5] ? way1_dirty_21 : _GEN_789; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_791 = 7'h16 == stage1_sram_addr_reg[11:5] ? way1_dirty_22 : _GEN_790; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_792 = 7'h17 == stage1_sram_addr_reg[11:5] ? way1_dirty_23 : _GEN_791; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_793 = 7'h18 == stage1_sram_addr_reg[11:5] ? way1_dirty_24 : _GEN_792; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_794 = 7'h19 == stage1_sram_addr_reg[11:5] ? way1_dirty_25 : _GEN_793; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_795 = 7'h1a == stage1_sram_addr_reg[11:5] ? way1_dirty_26 : _GEN_794; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_796 = 7'h1b == stage1_sram_addr_reg[11:5] ? way1_dirty_27 : _GEN_795; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_797 = 7'h1c == stage1_sram_addr_reg[11:5] ? way1_dirty_28 : _GEN_796; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_798 = 7'h1d == stage1_sram_addr_reg[11:5] ? way1_dirty_29 : _GEN_797; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_799 = 7'h1e == stage1_sram_addr_reg[11:5] ? way1_dirty_30 : _GEN_798; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_800 = 7'h1f == stage1_sram_addr_reg[11:5] ? way1_dirty_31 : _GEN_799; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_801 = 7'h20 == stage1_sram_addr_reg[11:5] ? way1_dirty_32 : _GEN_800; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_802 = 7'h21 == stage1_sram_addr_reg[11:5] ? way1_dirty_33 : _GEN_801; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_803 = 7'h22 == stage1_sram_addr_reg[11:5] ? way1_dirty_34 : _GEN_802; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_804 = 7'h23 == stage1_sram_addr_reg[11:5] ? way1_dirty_35 : _GEN_803; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_805 = 7'h24 == stage1_sram_addr_reg[11:5] ? way1_dirty_36 : _GEN_804; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_806 = 7'h25 == stage1_sram_addr_reg[11:5] ? way1_dirty_37 : _GEN_805; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_807 = 7'h26 == stage1_sram_addr_reg[11:5] ? way1_dirty_38 : _GEN_806; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_808 = 7'h27 == stage1_sram_addr_reg[11:5] ? way1_dirty_39 : _GEN_807; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_809 = 7'h28 == stage1_sram_addr_reg[11:5] ? way1_dirty_40 : _GEN_808; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_810 = 7'h29 == stage1_sram_addr_reg[11:5] ? way1_dirty_41 : _GEN_809; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_811 = 7'h2a == stage1_sram_addr_reg[11:5] ? way1_dirty_42 : _GEN_810; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_812 = 7'h2b == stage1_sram_addr_reg[11:5] ? way1_dirty_43 : _GEN_811; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_813 = 7'h2c == stage1_sram_addr_reg[11:5] ? way1_dirty_44 : _GEN_812; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_814 = 7'h2d == stage1_sram_addr_reg[11:5] ? way1_dirty_45 : _GEN_813; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_815 = 7'h2e == stage1_sram_addr_reg[11:5] ? way1_dirty_46 : _GEN_814; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_816 = 7'h2f == stage1_sram_addr_reg[11:5] ? way1_dirty_47 : _GEN_815; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_817 = 7'h30 == stage1_sram_addr_reg[11:5] ? way1_dirty_48 : _GEN_816; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_818 = 7'h31 == stage1_sram_addr_reg[11:5] ? way1_dirty_49 : _GEN_817; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_819 = 7'h32 == stage1_sram_addr_reg[11:5] ? way1_dirty_50 : _GEN_818; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_820 = 7'h33 == stage1_sram_addr_reg[11:5] ? way1_dirty_51 : _GEN_819; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_821 = 7'h34 == stage1_sram_addr_reg[11:5] ? way1_dirty_52 : _GEN_820; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_822 = 7'h35 == stage1_sram_addr_reg[11:5] ? way1_dirty_53 : _GEN_821; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_823 = 7'h36 == stage1_sram_addr_reg[11:5] ? way1_dirty_54 : _GEN_822; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_824 = 7'h37 == stage1_sram_addr_reg[11:5] ? way1_dirty_55 : _GEN_823; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_825 = 7'h38 == stage1_sram_addr_reg[11:5] ? way1_dirty_56 : _GEN_824; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_826 = 7'h39 == stage1_sram_addr_reg[11:5] ? way1_dirty_57 : _GEN_825; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_827 = 7'h3a == stage1_sram_addr_reg[11:5] ? way1_dirty_58 : _GEN_826; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_828 = 7'h3b == stage1_sram_addr_reg[11:5] ? way1_dirty_59 : _GEN_827; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_829 = 7'h3c == stage1_sram_addr_reg[11:5] ? way1_dirty_60 : _GEN_828; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_830 = 7'h3d == stage1_sram_addr_reg[11:5] ? way1_dirty_61 : _GEN_829; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_831 = 7'h3e == stage1_sram_addr_reg[11:5] ? way1_dirty_62 : _GEN_830; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_832 = 7'h3f == stage1_sram_addr_reg[11:5] ? way1_dirty_63 : _GEN_831; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_833 = 7'h40 == stage1_sram_addr_reg[11:5] ? way1_dirty_64 : _GEN_832; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_834 = 7'h41 == stage1_sram_addr_reg[11:5] ? way1_dirty_65 : _GEN_833; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_835 = 7'h42 == stage1_sram_addr_reg[11:5] ? way1_dirty_66 : _GEN_834; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_836 = 7'h43 == stage1_sram_addr_reg[11:5] ? way1_dirty_67 : _GEN_835; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_837 = 7'h44 == stage1_sram_addr_reg[11:5] ? way1_dirty_68 : _GEN_836; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_838 = 7'h45 == stage1_sram_addr_reg[11:5] ? way1_dirty_69 : _GEN_837; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_839 = 7'h46 == stage1_sram_addr_reg[11:5] ? way1_dirty_70 : _GEN_838; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_840 = 7'h47 == stage1_sram_addr_reg[11:5] ? way1_dirty_71 : _GEN_839; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_841 = 7'h48 == stage1_sram_addr_reg[11:5] ? way1_dirty_72 : _GEN_840; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_842 = 7'h49 == stage1_sram_addr_reg[11:5] ? way1_dirty_73 : _GEN_841; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_843 = 7'h4a == stage1_sram_addr_reg[11:5] ? way1_dirty_74 : _GEN_842; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_844 = 7'h4b == stage1_sram_addr_reg[11:5] ? way1_dirty_75 : _GEN_843; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_845 = 7'h4c == stage1_sram_addr_reg[11:5] ? way1_dirty_76 : _GEN_844; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_846 = 7'h4d == stage1_sram_addr_reg[11:5] ? way1_dirty_77 : _GEN_845; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_847 = 7'h4e == stage1_sram_addr_reg[11:5] ? way1_dirty_78 : _GEN_846; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_848 = 7'h4f == stage1_sram_addr_reg[11:5] ? way1_dirty_79 : _GEN_847; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_849 = 7'h50 == stage1_sram_addr_reg[11:5] ? way1_dirty_80 : _GEN_848; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_850 = 7'h51 == stage1_sram_addr_reg[11:5] ? way1_dirty_81 : _GEN_849; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_851 = 7'h52 == stage1_sram_addr_reg[11:5] ? way1_dirty_82 : _GEN_850; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_852 = 7'h53 == stage1_sram_addr_reg[11:5] ? way1_dirty_83 : _GEN_851; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_853 = 7'h54 == stage1_sram_addr_reg[11:5] ? way1_dirty_84 : _GEN_852; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_854 = 7'h55 == stage1_sram_addr_reg[11:5] ? way1_dirty_85 : _GEN_853; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_855 = 7'h56 == stage1_sram_addr_reg[11:5] ? way1_dirty_86 : _GEN_854; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_856 = 7'h57 == stage1_sram_addr_reg[11:5] ? way1_dirty_87 : _GEN_855; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_857 = 7'h58 == stage1_sram_addr_reg[11:5] ? way1_dirty_88 : _GEN_856; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_858 = 7'h59 == stage1_sram_addr_reg[11:5] ? way1_dirty_89 : _GEN_857; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_859 = 7'h5a == stage1_sram_addr_reg[11:5] ? way1_dirty_90 : _GEN_858; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_860 = 7'h5b == stage1_sram_addr_reg[11:5] ? way1_dirty_91 : _GEN_859; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_861 = 7'h5c == stage1_sram_addr_reg[11:5] ? way1_dirty_92 : _GEN_860; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_862 = 7'h5d == stage1_sram_addr_reg[11:5] ? way1_dirty_93 : _GEN_861; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_863 = 7'h5e == stage1_sram_addr_reg[11:5] ? way1_dirty_94 : _GEN_862; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_864 = 7'h5f == stage1_sram_addr_reg[11:5] ? way1_dirty_95 : _GEN_863; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_865 = 7'h60 == stage1_sram_addr_reg[11:5] ? way1_dirty_96 : _GEN_864; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_866 = 7'h61 == stage1_sram_addr_reg[11:5] ? way1_dirty_97 : _GEN_865; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_867 = 7'h62 == stage1_sram_addr_reg[11:5] ? way1_dirty_98 : _GEN_866; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_868 = 7'h63 == stage1_sram_addr_reg[11:5] ? way1_dirty_99 : _GEN_867; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_869 = 7'h64 == stage1_sram_addr_reg[11:5] ? way1_dirty_100 : _GEN_868; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_870 = 7'h65 == stage1_sram_addr_reg[11:5] ? way1_dirty_101 : _GEN_869; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_871 = 7'h66 == stage1_sram_addr_reg[11:5] ? way1_dirty_102 : _GEN_870; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_872 = 7'h67 == stage1_sram_addr_reg[11:5] ? way1_dirty_103 : _GEN_871; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_873 = 7'h68 == stage1_sram_addr_reg[11:5] ? way1_dirty_104 : _GEN_872; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_874 = 7'h69 == stage1_sram_addr_reg[11:5] ? way1_dirty_105 : _GEN_873; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_875 = 7'h6a == stage1_sram_addr_reg[11:5] ? way1_dirty_106 : _GEN_874; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_876 = 7'h6b == stage1_sram_addr_reg[11:5] ? way1_dirty_107 : _GEN_875; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_877 = 7'h6c == stage1_sram_addr_reg[11:5] ? way1_dirty_108 : _GEN_876; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_878 = 7'h6d == stage1_sram_addr_reg[11:5] ? way1_dirty_109 : _GEN_877; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_879 = 7'h6e == stage1_sram_addr_reg[11:5] ? way1_dirty_110 : _GEN_878; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_880 = 7'h6f == stage1_sram_addr_reg[11:5] ? way1_dirty_111 : _GEN_879; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_881 = 7'h70 == stage1_sram_addr_reg[11:5] ? way1_dirty_112 : _GEN_880; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_882 = 7'h71 == stage1_sram_addr_reg[11:5] ? way1_dirty_113 : _GEN_881; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_883 = 7'h72 == stage1_sram_addr_reg[11:5] ? way1_dirty_114 : _GEN_882; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_884 = 7'h73 == stage1_sram_addr_reg[11:5] ? way1_dirty_115 : _GEN_883; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_885 = 7'h74 == stage1_sram_addr_reg[11:5] ? way1_dirty_116 : _GEN_884; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_886 = 7'h75 == stage1_sram_addr_reg[11:5] ? way1_dirty_117 : _GEN_885; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_887 = 7'h76 == stage1_sram_addr_reg[11:5] ? way1_dirty_118 : _GEN_886; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_888 = 7'h77 == stage1_sram_addr_reg[11:5] ? way1_dirty_119 : _GEN_887; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_889 = 7'h78 == stage1_sram_addr_reg[11:5] ? way1_dirty_120 : _GEN_888; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_890 = 7'h79 == stage1_sram_addr_reg[11:5] ? way1_dirty_121 : _GEN_889; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_891 = 7'h7a == stage1_sram_addr_reg[11:5] ? way1_dirty_122 : _GEN_890; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_892 = 7'h7b == stage1_sram_addr_reg[11:5] ? way1_dirty_123 : _GEN_891; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_893 = 7'h7c == stage1_sram_addr_reg[11:5] ? way1_dirty_124 : _GEN_892; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_894 = 7'h7d == stage1_sram_addr_reg[11:5] ? way1_dirty_125 : _GEN_893; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_895 = 7'h7e == stage1_sram_addr_reg[11:5] ? way1_dirty_126 : _GEN_894; // @[data_cache.scala 157:{12,12}]
  wire  _GEN_896 = 7'h7f == stage1_sram_addr_reg[11:5] ? way1_dirty_127 : _GEN_895; // @[data_cache.scala 157:{12,12}]
  wire  _way1_dirty_T_14 = _way0_dirty_T_9 & _GEN_128 | _GEN_896; // @[data_cache.scala 157:12]
  wire  _way1_dirty_T_15 = _way0_dirty_T_5 & _GEN_128 ? 1'h0 : _way1_dirty_T_14; // @[data_cache.scala 156:12]
  wire  dirty_victim = _way0_dirty_T_7 ? _GEN_384 : _GEN_896; // @[data_cache.scala 161:24]
  wire  _io_tlb_req_T_4 = ~stage1_sram_addr_reg[31] | stage1_sram_addr_reg[31:30] == 2'h3; // @[macros.scala 424:18]
  wire [31:0] _stage1_sram_phy_addr_reg_T = io_tlb_req ? io_p_addr_for_tlb : stage1_sram_addr_reg; // @[data_cache.scala 176:73]
  wire [31:0] _stage1_sram_phy_addr_reg_T_4 = {3'h0,_stage1_sram_phy_addr_reg_T[28:0]}; // @[Cat.scala 31:58]
  wire  _lru_T_4 = _hit_T_1 ? 1'h0 : _GEN_128; // @[data_cache.scala 182:12]
  wire  _lru_T_5 = _hit_T | _lru_T_4; // @[data_cache.scala 181:12]
  wire [4:0] _state_ready_lookup_will_to_be_T_3 = stage1_sram_cache_reg ? 5'h19 : 5'h3; // @[data_cache.scala 190:16]
  wire [4:0] _state_ready_lookup_will_to_be_T_5 = stage1_sram_cache_reg ? 5'h19 : 5'h1; // @[data_cache.scala 190:88]
  wire [4:0] _state_ready_lookup_will_to_be_T_6 = stage1_sram_wr_reg ? _state_ready_lookup_will_to_be_T_3 :
    _state_ready_lookup_will_to_be_T_5; // @[data_cache.scala 189:81]
  wire [4:0] _state_ready_lookup_will_to_be_T_7 = stage1_sram_req_reg ? _state_ready_lookup_will_to_be_T_6 : 5'h19; // @[data_cache.scala 189:50]
  wire [1:0] _state_ready_lookup_will_to_be_T_12 = stage1_sram_wr_reg ? 2'h3 : 2'h1; // @[data_cache.scala 191:81]
  wire [3:0] _state_ready_lookup_will_to_be_T_15 = stage1_sram_wr_reg ? 4'h8 : 4'hc; // @[data_cache.scala 192:64]
  wire [3:0] _state_ready_lookup_will_to_be_T_16 = dirty_victim ? 4'h9 : _state_ready_lookup_will_to_be_T_15; // @[data_cache.scala 192:16]
  wire [3:0] _state_ready_lookup_will_to_be_T_17 = ~stage1_sram_cache_reg ? {{2'd0}, _state_ready_lookup_will_to_be_T_12
    } : _state_ready_lookup_will_to_be_T_16; // @[data_cache.scala 191:47]
  wire [4:0] _state_ready_lookup_will_to_be_T_18 = stage1_sram_req_reg ? {{1'd0}, _state_ready_lookup_will_to_be_T_17}
     : 5'h19; // @[data_cache.scala 191:16]
  wire [4:0] state_ready_lookup_will_to_be = hit ? _state_ready_lookup_will_to_be_T_7 :
    _state_ready_lookup_will_to_be_T_18; // @[data_cache.scala 189:42]
  wire [4:0] _access_work_state_T_1 = io_port_arready ? 5'h2 : work_state; // @[data_cache.scala 199:39]
  wire [4:0] _access_work_state_T_5 = io_port_awready ? 5'h4 : work_state; // @[data_cache.scala 202:39]
  wire [4:0] _access_work_state_T_7 = io_port_wready ? 5'h5 : work_state; // @[data_cache.scala 203:39]
  wire [4:0] _access_work_state_T_9 = io_port_arready ? 5'hd : work_state; // @[data_cache.scala 206:44]
  wire [4:0] _access_work_state_T_14 = stage1_sram_wr_reg ? 5'h10 : 5'he; // @[data_cache.scala 207:94]
  wire [4:0] _access_work_state_T_15 = io_port_rlast & io_port_rvalid ? _access_work_state_T_14 : work_state; // @[data_cache.scala 207:44]
  wire [4:0] _access_work_state_T_17 = io_port_awready ? 5'ha : work_state; // @[data_cache.scala 209:41]
  wire  _access_work_state_T_19 = write_counter == 3'h7; // @[data_cache.scala 210:81]
  wire  _access_work_state_T_20 = io_port_wready & write_counter == 3'h7; // @[data_cache.scala 210:64]
  wire [4:0] _access_work_state_T_21 = io_port_wready & write_counter == 3'h7 ? 5'hb : work_state; // @[data_cache.scala 210:41]
  wire [4:0] _access_work_state_T_23 = io_port_bvalid ? 5'hc : work_state; // @[data_cache.scala 211:41]
  wire [4:0] _access_work_state_T_25 = io_port_arready ? 5'h0 : work_state; // @[data_cache.scala 213:44]
  wire  _access_work_state_T_28 = io_port_rvalid & io_port_rlast; // @[data_cache.scala 214:68]
  wire [4:0] _access_work_state_T_29 = io_port_rvalid & io_port_rlast ? 5'h10 : work_state; // @[data_cache.scala 214:44]
  wire [4:0] _access_work_state_T_31 = io_port_awready ? 5'h6 : work_state; // @[data_cache.scala 216:41]
  wire [4:0] _access_work_state_T_39 = 5'h1 == work_state ? _access_work_state_T_1 : work_state; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_41 = 5'h2 == work_state ? _access_work_state_for_stall_T_1 : _access_work_state_T_39; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_43 = 5'h18 == work_state ? state_ready_lookup_will_to_be : _access_work_state_T_41; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_45 = 5'h3 == work_state ? _access_work_state_T_5 : _access_work_state_T_43; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_47 = 5'h4 == work_state ? _access_work_state_T_7 : _access_work_state_T_45; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_49 = 5'h5 == work_state ? 5'h18 : _access_work_state_T_47; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_51 = 5'h19 == work_state ? state_ready_lookup_will_to_be : _access_work_state_T_49; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_53 = 5'hc == work_state ? _access_work_state_T_9 : _access_work_state_T_51; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_55 = 5'hd == work_state ? _access_work_state_T_15 : _access_work_state_T_53; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_57 = 5'he == work_state ? 5'h18 : _access_work_state_T_55; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_59 = 5'h9 == work_state ? _access_work_state_T_17 : _access_work_state_T_57; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_61 = 5'ha == work_state ? _access_work_state_T_21 : _access_work_state_T_59; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_63 = 5'hb == work_state ? _access_work_state_T_23 : _access_work_state_T_61; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_65 = 5'h8 == work_state ? _access_work_state_T_25 : _access_work_state_T_63; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_67 = 5'h0 == work_state ? _access_work_state_T_29 : _access_work_state_T_65; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_69 = 5'h10 == work_state ? 5'h18 : _access_work_state_T_67; // @[Mux.scala 81:58]
  wire  _wait_data_T_3 = work_state == 5'hd; // @[data_cache.scala 237:24]
  wire  _write_counter_T = work_state == 5'ha; // @[data_cache.scala 239:37]
  wire [2:0] _write_counter_T_4 = write_counter + 3'h1; // @[data_cache.scala 239:139]
  wire [2:0] _write_counter_T_5 = _access_work_state_T_19 ? 3'h0 : _write_counter_T_4; // @[data_cache.scala 239:94]
  wire [2:0] _write_counter_T_6 = io_port_wready ? _write_counter_T_5 : write_counter; // @[data_cache.scala 239:68]
  wire  _write_counter_T_7 = work_state == 5'h6; // @[data_cache.scala 240:24]
  wire [2:0] _read_counter_T_6 = read_counter + 3'h1; // @[data_cache.scala 241:163]
  wire [2:0] _read_counter_T_7 = io_port_rvalid ? _read_counter_T_6 : read_counter; // @[data_cache.scala 241:128]
  wire [2:0] _read_counter_T_8 = _access_work_state_T_28 ? 3'h0 : _read_counter_T_7; // @[data_cache.scala 241:72]
  wire  _read_counter_T_9 = work_state == 5'h0; // @[data_cache.scala 242:24]
  reg [31:0] stage2_sram_addr_reg; // @[Reg.scala 28:20]
  reg  stage2_hit0_reg; // @[data_cache.scala 264:34]
  wire [31:0] dcache_data_way0_0_rdata = dcache_data_io_rdata; // @[data_cache.scala 70:{36,36}]
  wire [31:0] dcache_data_way0_1_rdata = dcache_data_1_io_rdata; // @[data_cache.scala 70:{36,36}]
  wire [31:0] _GEN_1923 = 3'h1 == stage2_sram_addr_reg[4:2] ? dcache_data_way0_1_rdata : dcache_data_way0_0_rdata; // @[data_cache.scala 289:{23,23}]
  wire [31:0] dcache_data_way0_2_rdata = dcache_data_2_io_rdata; // @[data_cache.scala 70:{36,36}]
  wire [31:0] _GEN_1924 = 3'h2 == stage2_sram_addr_reg[4:2] ? dcache_data_way0_2_rdata : _GEN_1923; // @[data_cache.scala 289:{23,23}]
  wire [31:0] dcache_data_way0_3_rdata = dcache_data_3_io_rdata; // @[data_cache.scala 70:{36,36}]
  wire [31:0] _GEN_1925 = 3'h3 == stage2_sram_addr_reg[4:2] ? dcache_data_way0_3_rdata : _GEN_1924; // @[data_cache.scala 289:{23,23}]
  wire [31:0] dcache_data_way0_4_rdata = dcache_data_4_io_rdata; // @[data_cache.scala 70:{36,36}]
  wire [31:0] _GEN_1926 = 3'h4 == stage2_sram_addr_reg[4:2] ? dcache_data_way0_4_rdata : _GEN_1925; // @[data_cache.scala 289:{23,23}]
  wire [31:0] dcache_data_way0_5_rdata = dcache_data_5_io_rdata; // @[data_cache.scala 70:{36,36}]
  wire [31:0] _GEN_1927 = 3'h5 == stage2_sram_addr_reg[4:2] ? dcache_data_way0_5_rdata : _GEN_1926; // @[data_cache.scala 289:{23,23}]
  wire [31:0] dcache_data_way0_6_rdata = dcache_data_6_io_rdata; // @[data_cache.scala 70:{36,36}]
  wire [31:0] _GEN_1928 = 3'h6 == stage2_sram_addr_reg[4:2] ? dcache_data_way0_6_rdata : _GEN_1927; // @[data_cache.scala 289:{23,23}]
  wire [31:0] dcache_data_way0_7_rdata = dcache_data_7_io_rdata; // @[data_cache.scala 70:{36,36}]
  wire [31:0] _GEN_1929 = 3'h7 == stage2_sram_addr_reg[4:2] ? dcache_data_way0_7_rdata : _GEN_1928; // @[data_cache.scala 289:{23,23}]
  wire [31:0] dcache_data_way1_0_rdata = dcache_data_8_io_rdata; // @[data_cache.scala 71:{36,36}]
  wire [31:0] dcache_data_way1_1_rdata = dcache_data_9_io_rdata; // @[data_cache.scala 71:{36,36}]
  wire [31:0] _GEN_1931 = 3'h1 == stage2_sram_addr_reg[4:2] ? dcache_data_way1_1_rdata : dcache_data_way1_0_rdata; // @[data_cache.scala 289:{23,23}]
  wire [31:0] dcache_data_way1_2_rdata = dcache_data_10_io_rdata; // @[data_cache.scala 71:{36,36}]
  wire [31:0] _GEN_1932 = 3'h2 == stage2_sram_addr_reg[4:2] ? dcache_data_way1_2_rdata : _GEN_1931; // @[data_cache.scala 289:{23,23}]
  wire [31:0] dcache_data_way1_3_rdata = dcache_data_11_io_rdata; // @[data_cache.scala 71:{36,36}]
  wire [31:0] _GEN_1933 = 3'h3 == stage2_sram_addr_reg[4:2] ? dcache_data_way1_3_rdata : _GEN_1932; // @[data_cache.scala 289:{23,23}]
  wire [31:0] dcache_data_way1_4_rdata = dcache_data_12_io_rdata; // @[data_cache.scala 71:{36,36}]
  wire [31:0] _GEN_1934 = 3'h4 == stage2_sram_addr_reg[4:2] ? dcache_data_way1_4_rdata : _GEN_1933; // @[data_cache.scala 289:{23,23}]
  wire [31:0] dcache_data_way1_5_rdata = dcache_data_13_io_rdata; // @[data_cache.scala 71:{36,36}]
  wire [31:0] _GEN_1935 = 3'h5 == stage2_sram_addr_reg[4:2] ? dcache_data_way1_5_rdata : _GEN_1934; // @[data_cache.scala 289:{23,23}]
  wire [31:0] dcache_data_way1_6_rdata = dcache_data_14_io_rdata; // @[data_cache.scala 71:{36,36}]
  wire [31:0] _GEN_1936 = 3'h6 == stage2_sram_addr_reg[4:2] ? dcache_data_way1_6_rdata : _GEN_1935; // @[data_cache.scala 289:{23,23}]
  wire [31:0] dcache_data_way1_7_rdata = dcache_data_15_io_rdata; // @[data_cache.scala 71:{36,36}]
  wire [31:0] _GEN_1937 = 3'h7 == stage2_sram_addr_reg[4:2] ? dcache_data_way1_7_rdata : _GEN_1936; // @[data_cache.scala 289:{23,23}]
  wire [31:0] hit_word = stage2_hit0_reg ? _GEN_1929 : _GEN_1937; // @[data_cache.scala 289:23]
  wire [31:0] _GEN_2067 = 3'h1 == write_counter ? dcache_data_way1_1_rdata : dcache_data_way1_0_rdata; // @[data_cache.scala 299:{29,29}]
  wire [31:0] _GEN_2068 = 3'h2 == write_counter ? dcache_data_way1_2_rdata : _GEN_2067; // @[data_cache.scala 299:{29,29}]
  wire [31:0] _GEN_2069 = 3'h3 == write_counter ? dcache_data_way1_3_rdata : _GEN_2068; // @[data_cache.scala 299:{29,29}]
  wire [31:0] _GEN_2070 = 3'h4 == write_counter ? dcache_data_way1_4_rdata : _GEN_2069; // @[data_cache.scala 299:{29,29}]
  wire [31:0] _GEN_2071 = 3'h5 == write_counter ? dcache_data_way1_5_rdata : _GEN_2070; // @[data_cache.scala 299:{29,29}]
  wire [31:0] _GEN_2072 = 3'h6 == write_counter ? dcache_data_way1_6_rdata : _GEN_2071; // @[data_cache.scala 299:{29,29}]
  wire [31:0] _GEN_2073 = 3'h7 == write_counter ? dcache_data_way1_7_rdata : _GEN_2072; // @[data_cache.scala 299:{29,29}]
  wire [31:0] _GEN_2075 = 3'h1 == write_counter ? dcache_data_way0_1_rdata : dcache_data_way0_0_rdata; // @[data_cache.scala 299:{29,29}]
  wire [31:0] _GEN_2076 = 3'h2 == write_counter ? dcache_data_way0_2_rdata : _GEN_2075; // @[data_cache.scala 299:{29,29}]
  wire [31:0] _GEN_2077 = 3'h3 == write_counter ? dcache_data_way0_3_rdata : _GEN_2076; // @[data_cache.scala 299:{29,29}]
  wire [31:0] _GEN_2078 = 3'h4 == write_counter ? dcache_data_way0_4_rdata : _GEN_2077; // @[data_cache.scala 299:{29,29}]
  wire [31:0] _GEN_2079 = 3'h5 == write_counter ? dcache_data_way0_5_rdata : _GEN_2078; // @[data_cache.scala 299:{29,29}]
  wire [31:0] _GEN_2080 = 3'h6 == write_counter ? dcache_data_way0_6_rdata : _GEN_2079; // @[data_cache.scala 299:{29,29}]
  wire [31:0] _GEN_2081 = 3'h7 == write_counter ? dcache_data_way0_7_rdata : _GEN_2080; // @[data_cache.scala 299:{29,29}]
  wire [31:0] writeback_data = _GEN_128 ? _GEN_2073 : _GEN_2081; // @[data_cache.scala 299:29]
  wire  _way0_burst_read_wen_T_2 = _wait_data_T_3 | _read_counter_T_9; // @[data_cache.scala 300:76]
  wire  _way0_burst_read_wen_T_4 = (_wait_data_T_3 | _read_counter_T_9) & io_port_rvalid; // @[data_cache.scala 300:124]
  wire  way0_burst_read_wen = (_wait_data_T_3 | _read_counter_T_9) & io_port_rvalid & _way0_dirty_T_7; // @[data_cache.scala 300:149]
  wire  way1_burst_read_wen = _way0_burst_read_wen_T_4 & _GEN_128; // @[data_cache.scala 301:149]
  wire  _dcache_data_way0_0_wdata_T_2 = _way0_dirty_T_9 | _way0_dirty_T; // @[data_cache.scala 304:81]
  wire [31:0] _dcache_data_way0_0_wdata_T_6 = _way0_burst_read_wen_T_2 ? io_port_rdata : 32'h0; // @[data_cache.scala 304:155]
  wire  _wen_way0_wire_0_T_1 = stage1_sram_addr_reg[4:2] == 3'h0; // @[data_cache.scala 314:61]
  wire  _way0_wen_0_T = 3'h0 == read_counter; // @[data_cache.scala 320:38]
  wire  way0_wen_0 = 3'h0 == read_counter & way0_burst_read_wen; // @[data_cache.scala 320:28]
  wire [3:0] _wen_way0_wire_0_T_13 = {way0_wen_0,way0_wen_0,way0_wen_0,way0_wen_0}; // @[Cat.scala 31:58]
  wire  way1_wen_0 = _way0_wen_0_T & way1_burst_read_wen; // @[data_cache.scala 321:28]
  wire [3:0] _wen_way1_wire_0_T_13 = {way1_wen_0,way1_wen_0,way1_wen_0,way1_wen_0}; // @[Cat.scala 31:58]
  wire  _wen_way0_wire_1_T_1 = stage1_sram_addr_reg[4:2] == 3'h1; // @[data_cache.scala 314:61]
  wire  _way0_wen_1_T = 3'h1 == read_counter; // @[data_cache.scala 320:38]
  wire  way0_wen_1 = 3'h1 == read_counter & way0_burst_read_wen; // @[data_cache.scala 320:28]
  wire [3:0] _wen_way0_wire_1_T_13 = {way0_wen_1,way0_wen_1,way0_wen_1,way0_wen_1}; // @[Cat.scala 31:58]
  wire  way1_wen_1 = _way0_wen_1_T & way1_burst_read_wen; // @[data_cache.scala 321:28]
  wire [3:0] _wen_way1_wire_1_T_13 = {way1_wen_1,way1_wen_1,way1_wen_1,way1_wen_1}; // @[Cat.scala 31:58]
  wire  _wen_way0_wire_2_T_1 = stage1_sram_addr_reg[4:2] == 3'h2; // @[data_cache.scala 314:61]
  wire  _way0_wen_2_T = 3'h2 == read_counter; // @[data_cache.scala 320:38]
  wire  way0_wen_2 = 3'h2 == read_counter & way0_burst_read_wen; // @[data_cache.scala 320:28]
  wire [3:0] _wen_way0_wire_2_T_13 = {way0_wen_2,way0_wen_2,way0_wen_2,way0_wen_2}; // @[Cat.scala 31:58]
  wire  way1_wen_2 = _way0_wen_2_T & way1_burst_read_wen; // @[data_cache.scala 321:28]
  wire [3:0] _wen_way1_wire_2_T_13 = {way1_wen_2,way1_wen_2,way1_wen_2,way1_wen_2}; // @[Cat.scala 31:58]
  wire  _wen_way0_wire_3_T_1 = stage1_sram_addr_reg[4:2] == 3'h3; // @[data_cache.scala 314:61]
  wire  _way0_wen_3_T = 3'h3 == read_counter; // @[data_cache.scala 320:38]
  wire  way0_wen_3 = 3'h3 == read_counter & way0_burst_read_wen; // @[data_cache.scala 320:28]
  wire [3:0] _wen_way0_wire_3_T_13 = {way0_wen_3,way0_wen_3,way0_wen_3,way0_wen_3}; // @[Cat.scala 31:58]
  wire  way1_wen_3 = _way0_wen_3_T & way1_burst_read_wen; // @[data_cache.scala 321:28]
  wire [3:0] _wen_way1_wire_3_T_13 = {way1_wen_3,way1_wen_3,way1_wen_3,way1_wen_3}; // @[Cat.scala 31:58]
  wire  _wen_way0_wire_4_T_1 = stage1_sram_addr_reg[4:2] == 3'h4; // @[data_cache.scala 314:61]
  wire  _way0_wen_4_T = 3'h4 == read_counter; // @[data_cache.scala 320:38]
  wire  way0_wen_4 = 3'h4 == read_counter & way0_burst_read_wen; // @[data_cache.scala 320:28]
  wire [3:0] _wen_way0_wire_4_T_13 = {way0_wen_4,way0_wen_4,way0_wen_4,way0_wen_4}; // @[Cat.scala 31:58]
  wire  way1_wen_4 = _way0_wen_4_T & way1_burst_read_wen; // @[data_cache.scala 321:28]
  wire [3:0] _wen_way1_wire_4_T_13 = {way1_wen_4,way1_wen_4,way1_wen_4,way1_wen_4}; // @[Cat.scala 31:58]
  wire  _wen_way0_wire_5_T_1 = stage1_sram_addr_reg[4:2] == 3'h5; // @[data_cache.scala 314:61]
  wire  _way0_wen_5_T = 3'h5 == read_counter; // @[data_cache.scala 320:38]
  wire  way0_wen_5 = 3'h5 == read_counter & way0_burst_read_wen; // @[data_cache.scala 320:28]
  wire [3:0] _wen_way0_wire_5_T_13 = {way0_wen_5,way0_wen_5,way0_wen_5,way0_wen_5}; // @[Cat.scala 31:58]
  wire  way1_wen_5 = _way0_wen_5_T & way1_burst_read_wen; // @[data_cache.scala 321:28]
  wire [3:0] _wen_way1_wire_5_T_13 = {way1_wen_5,way1_wen_5,way1_wen_5,way1_wen_5}; // @[Cat.scala 31:58]
  wire  _wen_way0_wire_6_T_1 = stage1_sram_addr_reg[4:2] == 3'h6; // @[data_cache.scala 314:61]
  wire  _way0_wen_6_T = 3'h6 == read_counter; // @[data_cache.scala 320:38]
  wire  way0_wen_6 = 3'h6 == read_counter & way0_burst_read_wen; // @[data_cache.scala 320:28]
  wire [3:0] _wen_way0_wire_6_T_13 = {way0_wen_6,way0_wen_6,way0_wen_6,way0_wen_6}; // @[Cat.scala 31:58]
  wire  way1_wen_6 = _way0_wen_6_T & way1_burst_read_wen; // @[data_cache.scala 321:28]
  wire [3:0] _wen_way1_wire_6_T_13 = {way1_wen_6,way1_wen_6,way1_wen_6,way1_wen_6}; // @[Cat.scala 31:58]
  wire  _wen_way0_wire_7_T_1 = stage1_sram_addr_reg[4:2] == 3'h7; // @[data_cache.scala 314:61]
  wire  _way0_wen_7_T = 3'h7 == read_counter; // @[data_cache.scala 320:38]
  wire  way0_wen_7 = 3'h7 == read_counter & way0_burst_read_wen; // @[data_cache.scala 320:28]
  wire [3:0] _wen_way0_wire_7_T_13 = {way0_wen_7,way0_wen_7,way0_wen_7,way0_wen_7}; // @[Cat.scala 31:58]
  wire  way1_wen_7 = _way0_wen_7_T & way1_burst_read_wen; // @[data_cache.scala 321:28]
  wire [3:0] _wen_way1_wire_7_T_13 = {way1_wen_7,way1_wen_7,way1_wen_7,way1_wen_7}; // @[Cat.scala 31:58]
  wire  _cache_wdata_T_3 = work_state == 5'h19; // @[data_cache.scala 327:24]
  wire [20:0] _T_21 = {1'h1,stage1_sram_addr_reg[31:12]}; // @[Cat.scala 31:58]
  wire  _io_port_araddr_T = work_state == 5'h1; // @[data_cache.scala 340:38]
  wire  _io_port_araddr_T_1 = work_state == 5'hc; // @[data_cache.scala 341:24]
  wire  _io_port_araddr_T_2 = work_state == 5'h8; // @[data_cache.scala 341:71]
  wire [31:0] _io_port_araddr_T_5 = {stage1_sram_phy_addr_reg[31:5],5'h0}; // @[Cat.scala 31:58]
  wire [31:0] _io_port_araddr_T_6 = work_state == 5'hc | work_state == 5'h8 ? _io_port_araddr_T_5 : 32'h0; // @[data_cache.scala 341:12]
  wire [2:0] _io_port_arlen_T_1 = stage1_sram_cache_reg ? 3'h7 : 3'h0; // @[data_cache.scala 342:26]
  wire [1:0] _io_port_arsize_T_1 = stage1_sram_cache_reg ? 2'h2 : stage1_sram_size_reg; // @[data_cache.scala 343:27]
  wire  stage2_addr_same_as_stage1 = stage2_sram_addr_reg == stage1_sram_addr_reg; // @[data_cache.scala 352:56]
  wire  stage2_write_stage1_read = stage2_sram_write_reg & ~stage1_sram_wr_reg; // @[data_cache.scala 353:58]
  wire  _T_29 = work_state == 5'h3; // @[data_cache.scala 354:21]
  wire  _GEN_4642 = io_port_bvalid ? 1'h0 : write_access_complete_reg; // @[data_cache.scala 356:39 357:35 359:35]
  wire [19:0] _awaddr_miss_addr_T_2 = _way0_dirty_T_7 ? dcache_tag_io_tag : dcache_tag_1_io_tag; // @[data_cache.scala 362:36]
  wire [31:0] awaddr_miss_addr = {_awaddr_miss_addr_T_2,stage1_sram_phy_addr_reg[11:5],5'h0}; // @[Cat.scala 31:58]
  wire  _io_port_arvalid_T_7 = ~(stage2_addr_same_as_stage1 & stage2_write_stage1_read & write_access_complete_reg); // @[data_cache.scala 365:53]
  wire  _io_port_arvalid_T_8 = (_io_port_araddr_T | _io_port_araddr_T_1 | _io_port_araddr_T_2) & _io_port_arvalid_T_7; // @[data_cache.scala 364:27]
  wire  _io_port_arvalid_T_10 = stage1_exception == 3'h0; // @[data_cache.scala 365:173]
  wire [31:0] _io_port_awaddr_T_2 = 5'h3 == work_state ? stage1_sram_phy_addr_reg : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_port_awaddr_T_4 = 5'h9 == work_state ? awaddr_miss_addr : _io_port_awaddr_T_2; // @[Mux.scala 81:58]
  wire  _io_port_wdata_T = work_state == 5'h4; // @[data_cache.scala 386:38]
  wire  _io_port_wdata_T_3 = _write_counter_T | _write_counter_T_7; // @[data_cache.scala 386:132]
  wire [31:0] _io_port_wdata_T_4 = _write_counter_T | _write_counter_T_7 ? writeback_data : 32'h0; // @[data_cache.scala 386:92]
  wire [3:0] _io_port_wstrb_T_4 = _io_port_wdata_T_3 ? 4'hf : 4'h0; // @[data_cache.scala 388:87]
  wire  _io_port_wlast_T_5 = _io_port_wdata_T_3 & _access_work_state_T_19; // @[data_cache.scala 391:9]
  wire  _io_port_sram_data_ok_T_1 = work_state == 5'h18; // @[data_cache.scala 397:79]
  reg [31:0] sram_rdata_reg; // @[data_cache.scala 398:33]
  reg  stage2_stall_reg; // @[data_cache.scala 400:35]
  wire [31:0] _io_port_sram_rdata_T_2 = _cache_wdata_T_3 ? hit_word : 32'h0; // @[data_cache.scala 402:97]
  wire [31:0] _io_port_sram_rdata_T_3 = _io_port_sram_data_ok_T_1 ? wait_data : _io_port_sram_rdata_T_2; // @[data_cache.scala 402:51]
  dcache_tag dcache_tag ( // @[data_cache.scala 37:30]
    .clock(dcache_tag_clock),
    .reset(dcache_tag_reset),
    .io_wen(dcache_tag_io_wen),
    .io_wdata(dcache_tag_io_wdata),
    .io_raddr(dcache_tag_io_raddr),
    .io_waddr(dcache_tag_io_waddr),
    .io_hit(dcache_tag_io_hit),
    .io_valid(dcache_tag_io_valid),
    .io_tag(dcache_tag_io_tag)
  );
  dcache_tag dcache_tag_1 ( // @[data_cache.scala 38:30]
    .clock(dcache_tag_1_clock),
    .reset(dcache_tag_1_reset),
    .io_wen(dcache_tag_1_io_wen),
    .io_wdata(dcache_tag_1_io_wdata),
    .io_raddr(dcache_tag_1_io_raddr),
    .io_waddr(dcache_tag_1_io_waddr),
    .io_hit(dcache_tag_1_io_hit),
    .io_valid(dcache_tag_1_io_valid),
    .io_tag(dcache_tag_1_io_tag)
  );
  dcache_data dcache_data ( // @[data_cache.scala 70:55]
    .clock(dcache_data_clock),
    .io_wen(dcache_data_io_wen),
    .io_addr(dcache_data_io_addr),
    .io_wdata(dcache_data_io_wdata),
    .io_rdata(dcache_data_io_rdata)
  );
  dcache_data dcache_data_1 ( // @[data_cache.scala 70:55]
    .clock(dcache_data_1_clock),
    .io_wen(dcache_data_1_io_wen),
    .io_addr(dcache_data_1_io_addr),
    .io_wdata(dcache_data_1_io_wdata),
    .io_rdata(dcache_data_1_io_rdata)
  );
  dcache_data dcache_data_2 ( // @[data_cache.scala 70:55]
    .clock(dcache_data_2_clock),
    .io_wen(dcache_data_2_io_wen),
    .io_addr(dcache_data_2_io_addr),
    .io_wdata(dcache_data_2_io_wdata),
    .io_rdata(dcache_data_2_io_rdata)
  );
  dcache_data dcache_data_3 ( // @[data_cache.scala 70:55]
    .clock(dcache_data_3_clock),
    .io_wen(dcache_data_3_io_wen),
    .io_addr(dcache_data_3_io_addr),
    .io_wdata(dcache_data_3_io_wdata),
    .io_rdata(dcache_data_3_io_rdata)
  );
  dcache_data dcache_data_4 ( // @[data_cache.scala 70:55]
    .clock(dcache_data_4_clock),
    .io_wen(dcache_data_4_io_wen),
    .io_addr(dcache_data_4_io_addr),
    .io_wdata(dcache_data_4_io_wdata),
    .io_rdata(dcache_data_4_io_rdata)
  );
  dcache_data dcache_data_5 ( // @[data_cache.scala 70:55]
    .clock(dcache_data_5_clock),
    .io_wen(dcache_data_5_io_wen),
    .io_addr(dcache_data_5_io_addr),
    .io_wdata(dcache_data_5_io_wdata),
    .io_rdata(dcache_data_5_io_rdata)
  );
  dcache_data dcache_data_6 ( // @[data_cache.scala 70:55]
    .clock(dcache_data_6_clock),
    .io_wen(dcache_data_6_io_wen),
    .io_addr(dcache_data_6_io_addr),
    .io_wdata(dcache_data_6_io_wdata),
    .io_rdata(dcache_data_6_io_rdata)
  );
  dcache_data dcache_data_7 ( // @[data_cache.scala 70:55]
    .clock(dcache_data_7_clock),
    .io_wen(dcache_data_7_io_wen),
    .io_addr(dcache_data_7_io_addr),
    .io_wdata(dcache_data_7_io_wdata),
    .io_rdata(dcache_data_7_io_rdata)
  );
  dcache_data dcache_data_8 ( // @[data_cache.scala 71:55]
    .clock(dcache_data_8_clock),
    .io_wen(dcache_data_8_io_wen),
    .io_addr(dcache_data_8_io_addr),
    .io_wdata(dcache_data_8_io_wdata),
    .io_rdata(dcache_data_8_io_rdata)
  );
  dcache_data dcache_data_9 ( // @[data_cache.scala 71:55]
    .clock(dcache_data_9_clock),
    .io_wen(dcache_data_9_io_wen),
    .io_addr(dcache_data_9_io_addr),
    .io_wdata(dcache_data_9_io_wdata),
    .io_rdata(dcache_data_9_io_rdata)
  );
  dcache_data dcache_data_10 ( // @[data_cache.scala 71:55]
    .clock(dcache_data_10_clock),
    .io_wen(dcache_data_10_io_wen),
    .io_addr(dcache_data_10_io_addr),
    .io_wdata(dcache_data_10_io_wdata),
    .io_rdata(dcache_data_10_io_rdata)
  );
  dcache_data dcache_data_11 ( // @[data_cache.scala 71:55]
    .clock(dcache_data_11_clock),
    .io_wen(dcache_data_11_io_wen),
    .io_addr(dcache_data_11_io_addr),
    .io_wdata(dcache_data_11_io_wdata),
    .io_rdata(dcache_data_11_io_rdata)
  );
  dcache_data dcache_data_12 ( // @[data_cache.scala 71:55]
    .clock(dcache_data_12_clock),
    .io_wen(dcache_data_12_io_wen),
    .io_addr(dcache_data_12_io_addr),
    .io_wdata(dcache_data_12_io_wdata),
    .io_rdata(dcache_data_12_io_rdata)
  );
  dcache_data dcache_data_13 ( // @[data_cache.scala 71:55]
    .clock(dcache_data_13_clock),
    .io_wen(dcache_data_13_io_wen),
    .io_addr(dcache_data_13_io_addr),
    .io_wdata(dcache_data_13_io_wdata),
    .io_rdata(dcache_data_13_io_rdata)
  );
  dcache_data dcache_data_14 ( // @[data_cache.scala 71:55]
    .clock(dcache_data_14_clock),
    .io_wen(dcache_data_14_io_wen),
    .io_addr(dcache_data_14_io_addr),
    .io_wdata(dcache_data_14_io_wdata),
    .io_rdata(dcache_data_14_io_rdata)
  );
  dcache_data dcache_data_15 ( // @[data_cache.scala 71:55]
    .clock(dcache_data_15_clock),
    .io_wen(dcache_data_15_io_wen),
    .io_addr(dcache_data_15_io_addr),
    .io_wdata(dcache_data_15_io_wdata),
    .io_rdata(dcache_data_15_io_rdata)
  );
  assign io_port_araddr = work_state == 5'h1 ? stage1_sram_phy_addr_reg : _io_port_araddr_T_6; // @[data_cache.scala 340:26]
  assign io_port_arlen = {{1'd0}, _io_port_arlen_T_1}; // @[data_cache.scala 342:20]
  assign io_port_arsize = {{1'd0}, _io_port_arsize_T_1}; // @[data_cache.scala 343:20]
  assign io_port_arburst = {{1'd0}, stage1_sram_cache_reg}; // @[data_cache.scala 347:21]
  assign io_port_arvalid = _io_port_arvalid_T_8 & stage1_exception == 3'h0; // @[data_cache.scala 365:153]
  assign io_port_awaddr = 5'hf == work_state ? awaddr_miss_addr : _io_port_awaddr_T_4; // @[Mux.scala 81:58]
  assign io_port_awlen = {{1'd0}, _io_port_arlen_T_1}; // @[data_cache.scala 374:21]
  assign io_port_awsize = {{1'd0}, _io_port_arsize_T_1}; // @[data_cache.scala 375:21]
  assign io_port_awburst = {{1'd0}, stage1_sram_cache_reg}; // @[data_cache.scala 379:21]
  assign io_port_awvalid = (_T_29 | work_state == 5'hf | work_state == 5'h9) & _io_port_arvalid_T_10; // @[data_cache.scala 383:168]
  assign io_port_wdata = work_state == 5'h4 ? stage1_sram_wdata_reg : _io_port_wdata_T_4; // @[data_cache.scala 386:26]
  assign io_port_wstrb = _io_port_wdata_T ? stage1_wstrb_reg : _io_port_wstrb_T_4; // @[data_cache.scala 388:26]
  assign io_port_wlast = _io_port_wdata_T | _io_port_wlast_T_5; // @[data_cache.scala 390:63]
  assign io_port_wvalid = _io_port_wdata_T | _write_counter_T | _write_counter_T_7; // @[data_cache.scala 392:105]
  assign io_port_sram_rdata = stage2_stall_reg ? _io_port_sram_rdata_T_3 : sram_rdata_reg; // @[data_cache.scala 402:30]
  assign io_stage2_stall = access_work_state_for_stall[4:3] == 2'h3 | stage1_exception != 3'h0; // @[data_cache.scala 232:66]
  assign io_stage1_wr = stage1_sram_wr_reg; // @[data_cache.scala 175:23]
  assign io_v_addr_for_tlb = stage1_sram_addr_reg; // @[data_cache.scala 174:23]
  assign io_tlb_req = _io_tlb_req_T_4 & stage1_sram_req_reg; // @[data_cache.scala 173:54]
  assign io_stage1_tlb_exception = stage1_exception; // @[data_cache.scala 276:29]
  assign dcache_tag_clock = clock;
  assign dcache_tag_reset = reset;
  assign dcache_tag_io_wen = _way0_burst_read_wen_T_2 & _way0_dirty_T_7; // @[data_cache.scala 330:122]
  assign dcache_tag_io_wdata = _way0_burst_read_wen_T_2 ? _T_21 : 21'h0; // @[data_cache.scala 332:30]
  assign dcache_tag_io_raddr = io_port_sram_addr; // @[data_cache.scala 168:24]
  assign dcache_tag_io_waddr = stage1_sram_addr_reg; // @[data_cache.scala 165:24]
  assign dcache_tag_1_clock = clock;
  assign dcache_tag_1_reset = reset;
  assign dcache_tag_1_io_wen = _way0_burst_read_wen_T_2 & _GEN_128; // @[data_cache.scala 331:122]
  assign dcache_tag_1_io_wdata = _way0_burst_read_wen_T_2 ? _T_21 : 21'h0; // @[data_cache.scala 333:30]
  assign dcache_tag_1_io_raddr = io_port_sram_addr; // @[data_cache.scala 169:24]
  assign dcache_tag_1_io_waddr = stage1_sram_addr_reg; // @[data_cache.scala 166:24]
  assign dcache_data_clock = clock;
  assign dcache_data_io_wen = stage1_sram_addr_reg[4:2] == 3'h0 & (_way0_dirty_T_4 | _way0_dirty_T_12) ?
    stage1_wstrb_reg : _wen_way0_wire_0_T_13; // @[data_cache.scala 314:33]
  assign dcache_data_io_addr = stage1_sram_addr_reg; // @[data_cache.scala 303:34 70:36]
  assign dcache_data_io_wdata = _way0_dirty_T_9 | _way0_dirty_T ? stage1_sram_wdata_reg : _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 304:41]
  assign dcache_data_1_clock = clock;
  assign dcache_data_1_io_wen = stage1_sram_addr_reg[4:2] == 3'h1 & (_way0_dirty_T_4 | _way0_dirty_T_12) ?
    stage1_wstrb_reg : _wen_way0_wire_1_T_13; // @[data_cache.scala 314:33]
  assign dcache_data_1_io_addr = stage1_sram_addr_reg; // @[data_cache.scala 303:34 70:36]
  assign dcache_data_1_io_wdata = _way0_dirty_T_9 | _way0_dirty_T ? stage1_sram_wdata_reg :
    _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 304:41]
  assign dcache_data_2_clock = clock;
  assign dcache_data_2_io_wen = stage1_sram_addr_reg[4:2] == 3'h2 & (_way0_dirty_T_4 | _way0_dirty_T_12) ?
    stage1_wstrb_reg : _wen_way0_wire_2_T_13; // @[data_cache.scala 314:33]
  assign dcache_data_2_io_addr = stage1_sram_addr_reg; // @[data_cache.scala 303:34 70:36]
  assign dcache_data_2_io_wdata = _way0_dirty_T_9 | _way0_dirty_T ? stage1_sram_wdata_reg :
    _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 304:41]
  assign dcache_data_3_clock = clock;
  assign dcache_data_3_io_wen = stage1_sram_addr_reg[4:2] == 3'h3 & (_way0_dirty_T_4 | _way0_dirty_T_12) ?
    stage1_wstrb_reg : _wen_way0_wire_3_T_13; // @[data_cache.scala 314:33]
  assign dcache_data_3_io_addr = stage1_sram_addr_reg; // @[data_cache.scala 303:34 70:36]
  assign dcache_data_3_io_wdata = _way0_dirty_T_9 | _way0_dirty_T ? stage1_sram_wdata_reg :
    _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 304:41]
  assign dcache_data_4_clock = clock;
  assign dcache_data_4_io_wen = stage1_sram_addr_reg[4:2] == 3'h4 & (_way0_dirty_T_4 | _way0_dirty_T_12) ?
    stage1_wstrb_reg : _wen_way0_wire_4_T_13; // @[data_cache.scala 314:33]
  assign dcache_data_4_io_addr = stage1_sram_addr_reg; // @[data_cache.scala 303:34 70:36]
  assign dcache_data_4_io_wdata = _way0_dirty_T_9 | _way0_dirty_T ? stage1_sram_wdata_reg :
    _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 304:41]
  assign dcache_data_5_clock = clock;
  assign dcache_data_5_io_wen = stage1_sram_addr_reg[4:2] == 3'h5 & (_way0_dirty_T_4 | _way0_dirty_T_12) ?
    stage1_wstrb_reg : _wen_way0_wire_5_T_13; // @[data_cache.scala 314:33]
  assign dcache_data_5_io_addr = stage1_sram_addr_reg; // @[data_cache.scala 303:34 70:36]
  assign dcache_data_5_io_wdata = _way0_dirty_T_9 | _way0_dirty_T ? stage1_sram_wdata_reg :
    _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 304:41]
  assign dcache_data_6_clock = clock;
  assign dcache_data_6_io_wen = stage1_sram_addr_reg[4:2] == 3'h6 & (_way0_dirty_T_4 | _way0_dirty_T_12) ?
    stage1_wstrb_reg : _wen_way0_wire_6_T_13; // @[data_cache.scala 314:33]
  assign dcache_data_6_io_addr = stage1_sram_addr_reg; // @[data_cache.scala 303:34 70:36]
  assign dcache_data_6_io_wdata = _way0_dirty_T_9 | _way0_dirty_T ? stage1_sram_wdata_reg :
    _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 304:41]
  assign dcache_data_7_clock = clock;
  assign dcache_data_7_io_wen = stage1_sram_addr_reg[4:2] == 3'h7 & (_way0_dirty_T_4 | _way0_dirty_T_12) ?
    stage1_wstrb_reg : _wen_way0_wire_7_T_13; // @[data_cache.scala 314:33]
  assign dcache_data_7_io_addr = stage1_sram_addr_reg; // @[data_cache.scala 303:34 70:36]
  assign dcache_data_7_io_wdata = _way0_dirty_T_9 | _way0_dirty_T ? stage1_sram_wdata_reg :
    _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 304:41]
  assign dcache_data_8_clock = clock;
  assign dcache_data_8_io_wen = _wen_way0_wire_0_T_1 & (_way1_dirty_T_4 | _way1_dirty_T_12) ? stage1_wstrb_reg :
    _wen_way1_wire_0_T_13; // @[data_cache.scala 316:33]
  assign dcache_data_8_io_addr = stage1_sram_addr_reg; // @[data_cache.scala 307:34 71:36]
  assign dcache_data_8_io_wdata = _dcache_data_way0_0_wdata_T_2 ? stage1_sram_wdata_reg : _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 308:41]
  assign dcache_data_9_clock = clock;
  assign dcache_data_9_io_wen = _wen_way0_wire_1_T_1 & (_way1_dirty_T_4 | _way1_dirty_T_12) ? stage1_wstrb_reg :
    _wen_way1_wire_1_T_13; // @[data_cache.scala 316:33]
  assign dcache_data_9_io_addr = stage1_sram_addr_reg; // @[data_cache.scala 307:34 71:36]
  assign dcache_data_9_io_wdata = _dcache_data_way0_0_wdata_T_2 ? stage1_sram_wdata_reg : _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 308:41]
  assign dcache_data_10_clock = clock;
  assign dcache_data_10_io_wen = _wen_way0_wire_2_T_1 & (_way1_dirty_T_4 | _way1_dirty_T_12) ? stage1_wstrb_reg :
    _wen_way1_wire_2_T_13; // @[data_cache.scala 316:33]
  assign dcache_data_10_io_addr = stage1_sram_addr_reg; // @[data_cache.scala 307:34 71:36]
  assign dcache_data_10_io_wdata = _dcache_data_way0_0_wdata_T_2 ? stage1_sram_wdata_reg : _dcache_data_way0_0_wdata_T_6
    ; // @[data_cache.scala 308:41]
  assign dcache_data_11_clock = clock;
  assign dcache_data_11_io_wen = _wen_way0_wire_3_T_1 & (_way1_dirty_T_4 | _way1_dirty_T_12) ? stage1_wstrb_reg :
    _wen_way1_wire_3_T_13; // @[data_cache.scala 316:33]
  assign dcache_data_11_io_addr = stage1_sram_addr_reg; // @[data_cache.scala 307:34 71:36]
  assign dcache_data_11_io_wdata = _dcache_data_way0_0_wdata_T_2 ? stage1_sram_wdata_reg : _dcache_data_way0_0_wdata_T_6
    ; // @[data_cache.scala 308:41]
  assign dcache_data_12_clock = clock;
  assign dcache_data_12_io_wen = _wen_way0_wire_4_T_1 & (_way1_dirty_T_4 | _way1_dirty_T_12) ? stage1_wstrb_reg :
    _wen_way1_wire_4_T_13; // @[data_cache.scala 316:33]
  assign dcache_data_12_io_addr = stage1_sram_addr_reg; // @[data_cache.scala 307:34 71:36]
  assign dcache_data_12_io_wdata = _dcache_data_way0_0_wdata_T_2 ? stage1_sram_wdata_reg : _dcache_data_way0_0_wdata_T_6
    ; // @[data_cache.scala 308:41]
  assign dcache_data_13_clock = clock;
  assign dcache_data_13_io_wen = _wen_way0_wire_5_T_1 & (_way1_dirty_T_4 | _way1_dirty_T_12) ? stage1_wstrb_reg :
    _wen_way1_wire_5_T_13; // @[data_cache.scala 316:33]
  assign dcache_data_13_io_addr = stage1_sram_addr_reg; // @[data_cache.scala 307:34 71:36]
  assign dcache_data_13_io_wdata = _dcache_data_way0_0_wdata_T_2 ? stage1_sram_wdata_reg : _dcache_data_way0_0_wdata_T_6
    ; // @[data_cache.scala 308:41]
  assign dcache_data_14_clock = clock;
  assign dcache_data_14_io_wen = _wen_way0_wire_6_T_1 & (_way1_dirty_T_4 | _way1_dirty_T_12) ? stage1_wstrb_reg :
    _wen_way1_wire_6_T_13; // @[data_cache.scala 316:33]
  assign dcache_data_14_io_addr = stage1_sram_addr_reg; // @[data_cache.scala 307:34 71:36]
  assign dcache_data_14_io_wdata = _dcache_data_way0_0_wdata_T_2 ? stage1_sram_wdata_reg : _dcache_data_way0_0_wdata_T_6
    ; // @[data_cache.scala 308:41]
  assign dcache_data_15_clock = clock;
  assign dcache_data_15_io_wen = _wen_way0_wire_7_T_1 & (_way1_dirty_T_4 | _way1_dirty_T_12) ? stage1_wstrb_reg :
    _wen_way1_wire_7_T_13; // @[data_cache.scala 316:33]
  assign dcache_data_15_io_addr = stage1_sram_addr_reg; // @[data_cache.scala 307:34 71:36]
  assign dcache_data_15_io_wdata = _dcache_data_way0_0_wdata_T_2 ? stage1_sram_wdata_reg : _dcache_data_way0_0_wdata_T_6
    ; // @[data_cache.scala 308:41]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 234:22]
      work_state <= 5'h18;
    end else if (_stage2_stall_T_2) begin // @[Mux.scala 81:58]
      work_state <= 5'h19; // @[data_cache.scala 218:41]
    end else if (5'h7 == work_state) begin // @[Mux.scala 81:58]
      if (io_port_bvalid) begin // @[data_cache.scala 217:41]
        work_state <= 5'h8;
      end
    end else if (5'h6 == work_state) begin // @[Mux.scala 81:58]
      if (_access_work_state_T_20) begin
        work_state <= 5'h7;
      end
    end else if (5'hf == work_state) begin
      work_state <= _access_work_state_T_31;
    end else begin
      work_state <= _access_work_state_T_69;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 239:25]
      write_counter <= 3'h0;
    end else if (work_state == 5'ha) begin // @[data_cache.scala 240:12]
      write_counter <= _write_counter_T_6;
    end else if (work_state == 5'h6) begin
      write_counter <= _write_counter_T_6;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 241:24]
      read_counter <= 3'h0;
    end else if (_wait_data_T_3) begin // @[data_cache.scala 242:12]
      read_counter <= _read_counter_T_8;
    end else if (work_state == 5'h0) begin
      read_counter <= _read_counter_T_8;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 236:21]
      wait_data <= 32'h0;
    end else if (work_state == 5'h2 & io_port_rvalid) begin // @[data_cache.scala 237:12]
      wait_data <= io_port_rdata;
    end else if (work_state == 5'hd & io_port_rvalid & read_counter == stage1_sram_addr_reg[4:2]) begin
      wait_data <= io_port_rdata;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_0 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h0 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_0 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_0 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_0 <= lru_127;
      end else begin
        lru_0 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_1 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h1 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_1 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_1 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_1 <= lru_127;
      end else begin
        lru_1 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_2 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h2 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_2 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_2 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_2 <= lru_127;
      end else begin
        lru_2 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_3 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h3 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_3 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_3 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_3 <= lru_127;
      end else begin
        lru_3 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_4 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h4 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_4 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_4 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_4 <= lru_127;
      end else begin
        lru_4 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_5 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h5 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_5 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_5 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_5 <= lru_127;
      end else begin
        lru_5 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_6 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h6 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_6 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_6 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_6 <= lru_127;
      end else begin
        lru_6 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_7 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h7 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_7 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_7 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_7 <= lru_127;
      end else begin
        lru_7 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_8 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h8 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_8 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_8 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_8 <= lru_127;
      end else begin
        lru_8 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_9 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h9 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_9 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_9 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_9 <= lru_127;
      end else begin
        lru_9 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_10 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'ha == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_10 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_10 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_10 <= lru_127;
      end else begin
        lru_10 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_11 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'hb == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_11 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_11 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_11 <= lru_127;
      end else begin
        lru_11 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_12 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'hc == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_12 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_12 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_12 <= lru_127;
      end else begin
        lru_12 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_13 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'hd == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_13 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_13 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_13 <= lru_127;
      end else begin
        lru_13 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_14 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'he == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_14 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_14 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_14 <= lru_127;
      end else begin
        lru_14 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_15 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'hf == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_15 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_15 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_15 <= lru_127;
      end else begin
        lru_15 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_16 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h10 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_16 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_16 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_16 <= lru_127;
      end else begin
        lru_16 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_17 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h11 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_17 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_17 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_17 <= lru_127;
      end else begin
        lru_17 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_18 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h12 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_18 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_18 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_18 <= lru_127;
      end else begin
        lru_18 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_19 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h13 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_19 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_19 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_19 <= lru_127;
      end else begin
        lru_19 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_20 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h14 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_20 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_20 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_20 <= lru_127;
      end else begin
        lru_20 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_21 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h15 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_21 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_21 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_21 <= lru_127;
      end else begin
        lru_21 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_22 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h16 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_22 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_22 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_22 <= lru_127;
      end else begin
        lru_22 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_23 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h17 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_23 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_23 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_23 <= lru_127;
      end else begin
        lru_23 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_24 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h18 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_24 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_24 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_24 <= lru_127;
      end else begin
        lru_24 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_25 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h19 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_25 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_25 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_25 <= lru_127;
      end else begin
        lru_25 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_26 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h1a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_26 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_26 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_26 <= lru_127;
      end else begin
        lru_26 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_27 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h1b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_27 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_27 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_27 <= lru_127;
      end else begin
        lru_27 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_28 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h1c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_28 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_28 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_28 <= lru_127;
      end else begin
        lru_28 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_29 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h1d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_29 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_29 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_29 <= lru_127;
      end else begin
        lru_29 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_30 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h1e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_30 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_30 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_30 <= lru_127;
      end else begin
        lru_30 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_31 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h1f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_31 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_31 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_31 <= lru_127;
      end else begin
        lru_31 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_32 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h20 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_32 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_32 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_32 <= lru_127;
      end else begin
        lru_32 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_33 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h21 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_33 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_33 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_33 <= lru_127;
      end else begin
        lru_33 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_34 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h22 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_34 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_34 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_34 <= lru_127;
      end else begin
        lru_34 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_35 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h23 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_35 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_35 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_35 <= lru_127;
      end else begin
        lru_35 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_36 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h24 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_36 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_36 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_36 <= lru_127;
      end else begin
        lru_36 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_37 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h25 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_37 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_37 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_37 <= lru_127;
      end else begin
        lru_37 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_38 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h26 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_38 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_38 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_38 <= lru_127;
      end else begin
        lru_38 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_39 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h27 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_39 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_39 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_39 <= lru_127;
      end else begin
        lru_39 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_40 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h28 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_40 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_40 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_40 <= lru_127;
      end else begin
        lru_40 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_41 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h29 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_41 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_41 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_41 <= lru_127;
      end else begin
        lru_41 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_42 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h2a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_42 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_42 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_42 <= lru_127;
      end else begin
        lru_42 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_43 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h2b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_43 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_43 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_43 <= lru_127;
      end else begin
        lru_43 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_44 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h2c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_44 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_44 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_44 <= lru_127;
      end else begin
        lru_44 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_45 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h2d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_45 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_45 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_45 <= lru_127;
      end else begin
        lru_45 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_46 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h2e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_46 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_46 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_46 <= lru_127;
      end else begin
        lru_46 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_47 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h2f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_47 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_47 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_47 <= lru_127;
      end else begin
        lru_47 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_48 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h30 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_48 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_48 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_48 <= lru_127;
      end else begin
        lru_48 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_49 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h31 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_49 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_49 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_49 <= lru_127;
      end else begin
        lru_49 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_50 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h32 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_50 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_50 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_50 <= lru_127;
      end else begin
        lru_50 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_51 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h33 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_51 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_51 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_51 <= lru_127;
      end else begin
        lru_51 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_52 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h34 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_52 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_52 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_52 <= lru_127;
      end else begin
        lru_52 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_53 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h35 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_53 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_53 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_53 <= lru_127;
      end else begin
        lru_53 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_54 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h36 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_54 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_54 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_54 <= lru_127;
      end else begin
        lru_54 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_55 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h37 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_55 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_55 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_55 <= lru_127;
      end else begin
        lru_55 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_56 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h38 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_56 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_56 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_56 <= lru_127;
      end else begin
        lru_56 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_57 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h39 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_57 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_57 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_57 <= lru_127;
      end else begin
        lru_57 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_58 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h3a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_58 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_58 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_58 <= lru_127;
      end else begin
        lru_58 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_59 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h3b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_59 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_59 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_59 <= lru_127;
      end else begin
        lru_59 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_60 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h3c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_60 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_60 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_60 <= lru_127;
      end else begin
        lru_60 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_61 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h3d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_61 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_61 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_61 <= lru_127;
      end else begin
        lru_61 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_62 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h3e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_62 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_62 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_62 <= lru_127;
      end else begin
        lru_62 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_63 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h3f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_63 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_63 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_63 <= lru_127;
      end else begin
        lru_63 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_64 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h40 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_64 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_64 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_64 <= lru_127;
      end else begin
        lru_64 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_65 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h41 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_65 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_65 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_65 <= lru_127;
      end else begin
        lru_65 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_66 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h42 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_66 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_66 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_66 <= lru_127;
      end else begin
        lru_66 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_67 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h43 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_67 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_67 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_67 <= lru_127;
      end else begin
        lru_67 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_68 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h44 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_68 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_68 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_68 <= lru_127;
      end else begin
        lru_68 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_69 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h45 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_69 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_69 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_69 <= lru_127;
      end else begin
        lru_69 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_70 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h46 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_70 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_70 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_70 <= lru_127;
      end else begin
        lru_70 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_71 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h47 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_71 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_71 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_71 <= lru_127;
      end else begin
        lru_71 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_72 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h48 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_72 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_72 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_72 <= lru_127;
      end else begin
        lru_72 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_73 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h49 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_73 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_73 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_73 <= lru_127;
      end else begin
        lru_73 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_74 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h4a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_74 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_74 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_74 <= lru_127;
      end else begin
        lru_74 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_75 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h4b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_75 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_75 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_75 <= lru_127;
      end else begin
        lru_75 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_76 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h4c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_76 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_76 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_76 <= lru_127;
      end else begin
        lru_76 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_77 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h4d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_77 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_77 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_77 <= lru_127;
      end else begin
        lru_77 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_78 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h4e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_78 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_78 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_78 <= lru_127;
      end else begin
        lru_78 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_79 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h4f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_79 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_79 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_79 <= lru_127;
      end else begin
        lru_79 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_80 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h50 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_80 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_80 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_80 <= lru_127;
      end else begin
        lru_80 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_81 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h51 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_81 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_81 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_81 <= lru_127;
      end else begin
        lru_81 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_82 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h52 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_82 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_82 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_82 <= lru_127;
      end else begin
        lru_82 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_83 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h53 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_83 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_83 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_83 <= lru_127;
      end else begin
        lru_83 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_84 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h54 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_84 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_84 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_84 <= lru_127;
      end else begin
        lru_84 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_85 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h55 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_85 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_85 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_85 <= lru_127;
      end else begin
        lru_85 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_86 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h56 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_86 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_86 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_86 <= lru_127;
      end else begin
        lru_86 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_87 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h57 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_87 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_87 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_87 <= lru_127;
      end else begin
        lru_87 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_88 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h58 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_88 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_88 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_88 <= lru_127;
      end else begin
        lru_88 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_89 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h59 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_89 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_89 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_89 <= lru_127;
      end else begin
        lru_89 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_90 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h5a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_90 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_90 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_90 <= lru_127;
      end else begin
        lru_90 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_91 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h5b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_91 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_91 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_91 <= lru_127;
      end else begin
        lru_91 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_92 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h5c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_92 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_92 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_92 <= lru_127;
      end else begin
        lru_92 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_93 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h5d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_93 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_93 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_93 <= lru_127;
      end else begin
        lru_93 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_94 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h5e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_94 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_94 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_94 <= lru_127;
      end else begin
        lru_94 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_95 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h5f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_95 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_95 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_95 <= lru_127;
      end else begin
        lru_95 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_96 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h60 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_96 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_96 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_96 <= lru_127;
      end else begin
        lru_96 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_97 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h61 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_97 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_97 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_97 <= lru_127;
      end else begin
        lru_97 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_98 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h62 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_98 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_98 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_98 <= lru_127;
      end else begin
        lru_98 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_99 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h63 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_99 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_99 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_99 <= lru_127;
      end else begin
        lru_99 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_100 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h64 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_100 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_100 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_100 <= lru_127;
      end else begin
        lru_100 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_101 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h65 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_101 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_101 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_101 <= lru_127;
      end else begin
        lru_101 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_102 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h66 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_102 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_102 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_102 <= lru_127;
      end else begin
        lru_102 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_103 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h67 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_103 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_103 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_103 <= lru_127;
      end else begin
        lru_103 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_104 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h68 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_104 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_104 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_104 <= lru_127;
      end else begin
        lru_104 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_105 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h69 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_105 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_105 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_105 <= lru_127;
      end else begin
        lru_105 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_106 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h6a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_106 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_106 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_106 <= lru_127;
      end else begin
        lru_106 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_107 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h6b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_107 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_107 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_107 <= lru_127;
      end else begin
        lru_107 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_108 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h6c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_108 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_108 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_108 <= lru_127;
      end else begin
        lru_108 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_109 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h6d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_109 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_109 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_109 <= lru_127;
      end else begin
        lru_109 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_110 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h6e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_110 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_110 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_110 <= lru_127;
      end else begin
        lru_110 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_111 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h6f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_111 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_111 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_111 <= lru_127;
      end else begin
        lru_111 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_112 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h70 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_112 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_112 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_112 <= lru_127;
      end else begin
        lru_112 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_113 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h71 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_113 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_113 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_113 <= lru_127;
      end else begin
        lru_113 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_114 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h72 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_114 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_114 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_114 <= lru_127;
      end else begin
        lru_114 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_115 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h73 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_115 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_115 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_115 <= lru_127;
      end else begin
        lru_115 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_116 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h74 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_116 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_116 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_116 <= lru_127;
      end else begin
        lru_116 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_117 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h75 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_117 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_117 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_117 <= lru_127;
      end else begin
        lru_117 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_118 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h76 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_118 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_118 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_118 <= lru_127;
      end else begin
        lru_118 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_119 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h77 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_119 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_119 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_119 <= lru_127;
      end else begin
        lru_119 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_120 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h78 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_120 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_120 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_120 <= lru_127;
      end else begin
        lru_120 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_121 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h79 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_121 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_121 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_121 <= lru_127;
      end else begin
        lru_121 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_122 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h7a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_122 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_122 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_122 <= lru_127;
      end else begin
        lru_122 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_123 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h7b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_123 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_123 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_123 <= lru_127;
      end else begin
        lru_123 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_124 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h7c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_124 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_124 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_124 <= lru_127;
      end else begin
        lru_124 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_125 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h7d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_125 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_125 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_125 <= lru_127;
      end else begin
        lru_125 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_126 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h7e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_126 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_126 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin
        lru_126 <= lru_127;
      end else begin
        lru_126 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 180:37]
      lru_127 <= 1'h0; // @[data_cache.scala 180:43 183:12 152:{86,86}]
    end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 40:22]
      if (_way0_dirty_T) begin
        lru_127 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_127 <= _way0_dirty_T_7;
      end else if (!(7'h7f == stage1_sram_addr_reg[11:5])) begin
        lru_127 <= _GEN_127;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_0 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h0 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_0 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_1 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h1 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_1 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_2 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h2 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_2 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_3 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h3 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_3 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_4 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h4 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_4 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_5 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h5 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_5 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_6 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h6 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_6 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_7 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h7 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_7 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_8 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h8 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_8 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_9 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h9 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_9 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_10 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'ha == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_10 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_11 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'hb == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_11 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_12 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'hc == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_12 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_13 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'hd == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_13 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_14 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'he == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_14 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_15 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'hf == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_15 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_16 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h10 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_16 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_17 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h11 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_17 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_18 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h12 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_18 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_19 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h13 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_19 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_20 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h14 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_20 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_21 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h15 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_21 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_22 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h16 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_22 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_23 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h17 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_23 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_24 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h18 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_24 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_25 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h19 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_25 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_26 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h1a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_26 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_27 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h1b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_27 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_28 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h1c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_28 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_29 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h1d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_29 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_30 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h1e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_30 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_31 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h1f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_31 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_32 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h20 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_32 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_33 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h21 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_33 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_34 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h22 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_34 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_35 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h23 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_35 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_36 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h24 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_36 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_37 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h25 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_37 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_38 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h26 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_38 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_39 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h27 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_39 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_40 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h28 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_40 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_41 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h29 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_41 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_42 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h2a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_42 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_43 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h2b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_43 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_44 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h2c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_44 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_45 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h2d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_45 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_46 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h2e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_46 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_47 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h2f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_47 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_48 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h30 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_48 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_49 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h31 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_49 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_50 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h32 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_50 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_51 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h33 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_51 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_52 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h34 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_52 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_53 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h35 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_53 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_54 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h36 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_54 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_55 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h37 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_55 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_56 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h38 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_56 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_57 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h39 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_57 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_58 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h3a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_58 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_59 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h3b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_59 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_60 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h3c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_60 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_61 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h3d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_61 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_62 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h3e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_62 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_63 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h3f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_63 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_64 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h40 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_64 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_65 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h41 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_65 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_66 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h42 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_66 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_67 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h43 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_67 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_68 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h44 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_68 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_69 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h45 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_69 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_70 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h46 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_70 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_71 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h47 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_71 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_72 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h48 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_72 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_73 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h49 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_73 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_74 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h4a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_74 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_75 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h4b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_75 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_76 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h4c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_76 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_77 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h4d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_77 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_78 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h4e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_78 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_79 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h4f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_79 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_80 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h50 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_80 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_81 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h51 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_81 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_82 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h52 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_82 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_83 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h53 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_83 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_84 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h54 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_84 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_85 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h55 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_85 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_86 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h56 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_86 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_87 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h57 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_87 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_88 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h58 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_88 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_89 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h59 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_89 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_90 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h5a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_90 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_91 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h5b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_91 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_92 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h5c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_92 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_93 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h5d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_93 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_94 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h5e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_94 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_95 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h5f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_95 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_96 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h60 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_96 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_97 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h61 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_97 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_98 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h62 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_98 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_99 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h63 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_99 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_100 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h64 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_100 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_101 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h65 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_101 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_102 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h66 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_102 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_103 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h67 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_103 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_104 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h68 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_104 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_105 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h69 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_105 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_106 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h6a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_106 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_107 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h6b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_107 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_108 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h6c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_108 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_109 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h6d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_109 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_110 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h6e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_110 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_111 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h6f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_111 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_112 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h70 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_112 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_113 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h71 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_113 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_114 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h72 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_114 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_115 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h73 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_115 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_116 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h74 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_116 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_117 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h75 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_117 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_118 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h76 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_118 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_119 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h77 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_119 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_120 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h78 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_120 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_121 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h79 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_121 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_122 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h7a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_122 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_123 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h7b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_123 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_124 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h7c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_124 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_125 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h7d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_125 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_126 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h7e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_126 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 151:44]
      way0_dirty_127 <= 1'h0; // @[data_cache.scala 151:44]
    end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 41:29]
      way0_dirty_127 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_0 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h0 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_0 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_1 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h1 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_1 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_2 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h2 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_2 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_3 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h3 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_3 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_4 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h4 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_4 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_5 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h5 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_5 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_6 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h6 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_6 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_7 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h7 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_7 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_8 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h8 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_8 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_9 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h9 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_9 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_10 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'ha == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_10 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_11 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'hb == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_11 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_12 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'hc == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_12 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_13 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'hd == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_13 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_14 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'he == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_14 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_15 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'hf == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_15 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_16 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h10 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_16 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_17 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h11 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_17 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_18 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h12 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_18 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_19 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h13 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_19 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_20 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h14 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_20 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_21 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h15 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_21 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_22 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h16 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_22 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_23 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h17 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_23 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_24 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h18 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_24 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_25 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h19 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_25 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_26 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h1a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_26 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_27 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h1b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_27 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_28 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h1c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_28 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_29 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h1d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_29 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_30 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h1e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_30 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_31 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h1f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_31 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_32 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h20 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_32 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_33 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h21 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_33 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_34 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h22 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_34 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_35 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h23 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_35 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_36 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h24 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_36 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_37 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h25 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_37 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_38 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h26 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_38 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_39 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h27 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_39 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_40 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h28 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_40 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_41 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h29 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_41 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_42 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h2a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_42 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_43 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h2b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_43 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_44 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h2c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_44 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_45 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h2d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_45 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_46 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h2e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_46 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_47 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h2f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_47 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_48 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h30 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_48 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_49 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h31 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_49 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_50 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h32 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_50 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_51 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h33 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_51 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_52 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h34 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_52 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_53 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h35 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_53 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_54 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h36 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_54 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_55 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h37 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_55 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_56 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h38 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_56 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_57 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h39 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_57 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_58 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h3a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_58 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_59 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h3b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_59 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_60 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h3c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_60 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_61 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h3d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_61 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_62 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h3e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_62 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_63 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h3f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_63 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_64 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h40 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_64 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_65 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h41 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_65 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_66 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h42 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_66 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_67 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h43 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_67 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_68 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h44 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_68 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_69 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h45 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_69 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_70 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h46 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_70 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_71 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h47 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_71 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_72 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h48 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_72 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_73 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h49 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_73 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_74 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h4a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_74 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_75 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h4b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_75 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_76 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h4c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_76 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_77 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h4d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_77 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_78 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h4e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_78 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_79 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h4f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_79 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_80 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h50 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_80 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_81 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h51 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_81 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_82 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h52 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_82 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_83 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h53 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_83 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_84 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h54 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_84 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_85 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h55 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_85 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_86 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h56 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_86 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_87 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h57 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_87 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_88 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h58 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_88 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_89 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h59 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_89 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_90 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h5a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_90 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_91 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h5b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_91 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_92 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h5c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_92 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_93 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h5d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_93 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_94 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h5e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_94 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_95 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h5f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_95 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_96 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h60 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_96 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_97 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h61 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_97 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_98 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h62 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_98 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_99 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h63 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_99 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_100 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h64 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_100 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_101 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h65 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_101 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_102 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h66 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_102 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_103 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h67 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_103 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_104 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h68 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_104 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_105 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h69 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_105 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_106 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h6a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_106 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_107 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h6b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_107 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_108 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h6c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_108 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_109 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h6d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_109 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_110 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h6e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_110 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_111 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h6f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_111 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_112 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h70 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_112 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_113 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h71 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_113 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_114 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h72 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_114 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_115 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h73 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_115 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_116 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h74 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_116 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_117 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h75 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_117 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_118 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h76 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_118 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_119 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h77 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_119 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_120 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h78 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_120 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_121 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h79 == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_121 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_122 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h7a == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_122 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_123 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h7b == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_123 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_124 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h7c == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_124 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_125 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h7d == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_125 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_126 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h7e == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_126 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 155:44]
      way1_dirty_127 <= 1'h0; // @[data_cache.scala 155:44]
    end else if (7'h7f == stage1_sram_addr_reg[11:5]) begin // @[data_cache.scala 42:29]
      way1_dirty_127 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 137:32]
      stage1_sram_addr_reg <= 32'h0;
    end else if (io_port_sram_req) begin
      stage1_sram_addr_reg <= io_port_sram_addr;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 138:33]
      stage1_sram_cache_reg <= 1'h0;
    end else if (io_port_sram_req) begin
      stage1_sram_cache_reg <= io_port_sram_cache;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 139:33]
      stage1_sram_wdata_reg <= 32'h0;
    end else if (io_port_sram_req) begin
      stage1_sram_wdata_reg <= io_port_sram_wdata;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 140:33]
      stage1_sram_size_reg <= 2'h0;
    end else if (io_port_sram_req) begin
      stage1_sram_size_reg <= io_port_sram_size;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 141:33]
      stage1_sram_wr_reg <= 1'h0;
    end else if (io_port_sram_req) begin
      stage1_sram_wr_reg <= io_port_sram_wr;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 142:33]
      stage1_sram_req_reg <= 1'h0;
    end else begin
      stage1_sram_req_reg <= io_port_sram_req | _stage1_sram_req_reg_T_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 145:32]
      stage1_sram_hit0_reg <= 1'h0;
    end else if (io_port_sram_req) begin
      stage1_sram_hit0_reg <= dcache_tag_io_hit;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 146:32]
      stage1_sram_hit1_reg <= 1'h0;
    end else if (io_port_sram_req) begin
      stage1_sram_hit1_reg <= dcache_tag_1_io_hit;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 147:34]
      stage1_sram_valid0_reg <= 1'h0;
    end else if (io_port_sram_req) begin
      stage1_sram_valid0_reg <= dcache_tag_io_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 148:34]
      stage1_sram_valid1_reg <= 1'h0;
    end else if (io_port_sram_req) begin
      stage1_sram_valid1_reg <= dcache_tag_1_io_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 143:33]
      stage1_wstrb_reg <= 4'h0;
    end else if (io_port_sram_req) begin
      stage1_wstrb_reg <= io_data_wstrb;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 176:37]
      stage1_sram_phy_addr_reg <= 32'h0; // @[macros.scala 421:45 data_cache.scala 176:73]
    end else if (stage1_stall_reg) begin
      if (_stage1_sram_phy_addr_reg_T[31:30] == 2'h2) begin
        stage1_sram_phy_addr_reg <= _stage1_sram_phy_addr_reg_T_4;
      end else if (io_tlb_req) begin
        stage1_sram_phy_addr_reg <= io_p_addr_for_tlb;
      end else begin
        stage1_sram_phy_addr_reg <= stage1_sram_addr_reg;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 177:28]
      stage1_exception <= 3'h0;
    end else if (stage2_stall) begin
      stage1_exception <= 3'h0;
    end else begin
      stage1_exception <= io_tlb_exception;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 261:54]
      stage2_sram_write_reg <= 1'h0;
    end else if (stage2_stall) begin
      stage2_sram_write_reg <= stage1_sram_wr_reg;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 131:42]
      stage1_stall_reg <= 1'h0;
    end else begin
      stage1_stall_reg <= io_port_sram_req;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 354:52]
      write_access_complete_reg <= 1'h0; // @[data_cache.scala 355:35]
    end else begin
      write_access_complete_reg <= work_state == 5'h3 | _GEN_4642;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      stage2_sram_addr_reg <= 32'h0; // @[Reg.scala 29:22]
    end else if (stage2_stall) begin // @[Reg.scala 28:20]
      stage2_sram_addr_reg <= stage1_sram_addr_reg;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 265:48]
      stage2_hit0_reg <= 1'h0;
    end else if (stage2_stall) begin
      stage2_hit0_reg <= _hit_T;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 399:27]
      sram_rdata_reg <= 32'h0;
    end else if (_io_port_sram_data_ok_T_1) begin // @[data_cache.scala 399:73]
      sram_rdata_reg <= wait_data; // @[data_cache.scala 289:{23,23,23,23,23}]
    end else if (_cache_wdata_T_3) begin
      if (stage2_hit0_reg) begin
        if (3'h7 == stage2_sram_addr_reg[4:2]) begin
          sram_rdata_reg <= dcache_data_way0_7_rdata;
        end else begin
          sram_rdata_reg <= _GEN_1928;
        end
      end else if (3'h7 == stage2_sram_addr_reg[4:2]) begin
        sram_rdata_reg <= dcache_data_way1_7_rdata;
      end else begin
        sram_rdata_reg <= _GEN_1936;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 232:66]
      stage2_stall_reg <= 1'h0;
    end else begin
      stage2_stall_reg <= access_work_state_for_stall[4:3] == 2'h3 | stage1_exception != 3'h0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  work_state = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  write_counter = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  read_counter = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  wait_data = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  lru_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lru_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  lru_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  lru_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  lru_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  lru_5 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  lru_6 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  lru_7 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  lru_8 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  lru_9 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  lru_10 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  lru_11 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  lru_12 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  lru_13 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  lru_14 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  lru_15 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  lru_16 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  lru_17 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  lru_18 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  lru_19 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  lru_20 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  lru_21 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  lru_22 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  lru_23 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  lru_24 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  lru_25 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  lru_26 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  lru_27 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  lru_28 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  lru_29 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  lru_30 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  lru_31 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  lru_32 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  lru_33 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  lru_34 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  lru_35 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  lru_36 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  lru_37 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  lru_38 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  lru_39 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  lru_40 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  lru_41 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  lru_42 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  lru_43 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  lru_44 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  lru_45 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  lru_46 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  lru_47 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  lru_48 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  lru_49 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  lru_50 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  lru_51 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  lru_52 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  lru_53 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  lru_54 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  lru_55 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  lru_56 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  lru_57 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  lru_58 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  lru_59 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  lru_60 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  lru_61 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  lru_62 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  lru_63 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  lru_64 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  lru_65 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  lru_66 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  lru_67 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  lru_68 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  lru_69 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  lru_70 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  lru_71 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  lru_72 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  lru_73 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  lru_74 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  lru_75 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  lru_76 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  lru_77 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  lru_78 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  lru_79 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  lru_80 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  lru_81 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  lru_82 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  lru_83 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  lru_84 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  lru_85 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  lru_86 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  lru_87 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  lru_88 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  lru_89 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  lru_90 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  lru_91 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  lru_92 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  lru_93 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  lru_94 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  lru_95 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  lru_96 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  lru_97 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  lru_98 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  lru_99 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  lru_100 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  lru_101 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  lru_102 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  lru_103 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  lru_104 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  lru_105 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  lru_106 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  lru_107 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  lru_108 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  lru_109 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  lru_110 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  lru_111 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  lru_112 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  lru_113 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  lru_114 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  lru_115 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  lru_116 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  lru_117 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  lru_118 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  lru_119 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  lru_120 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  lru_121 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  lru_122 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  lru_123 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  lru_124 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  lru_125 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  lru_126 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  lru_127 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  way0_dirty_0 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  way0_dirty_1 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  way0_dirty_2 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  way0_dirty_3 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  way0_dirty_4 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  way0_dirty_5 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  way0_dirty_6 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  way0_dirty_7 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  way0_dirty_8 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  way0_dirty_9 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  way0_dirty_10 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  way0_dirty_11 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  way0_dirty_12 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  way0_dirty_13 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  way0_dirty_14 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  way0_dirty_15 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  way0_dirty_16 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  way0_dirty_17 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  way0_dirty_18 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  way0_dirty_19 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  way0_dirty_20 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  way0_dirty_21 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  way0_dirty_22 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  way0_dirty_23 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  way0_dirty_24 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  way0_dirty_25 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  way0_dirty_26 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  way0_dirty_27 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  way0_dirty_28 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  way0_dirty_29 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  way0_dirty_30 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  way0_dirty_31 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  way0_dirty_32 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  way0_dirty_33 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  way0_dirty_34 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  way0_dirty_35 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  way0_dirty_36 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  way0_dirty_37 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  way0_dirty_38 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  way0_dirty_39 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  way0_dirty_40 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  way0_dirty_41 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  way0_dirty_42 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  way0_dirty_43 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  way0_dirty_44 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  way0_dirty_45 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  way0_dirty_46 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  way0_dirty_47 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  way0_dirty_48 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  way0_dirty_49 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  way0_dirty_50 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  way0_dirty_51 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  way0_dirty_52 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  way0_dirty_53 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  way0_dirty_54 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  way0_dirty_55 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  way0_dirty_56 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  way0_dirty_57 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  way0_dirty_58 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  way0_dirty_59 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  way0_dirty_60 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  way0_dirty_61 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  way0_dirty_62 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  way0_dirty_63 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  way0_dirty_64 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  way0_dirty_65 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  way0_dirty_66 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  way0_dirty_67 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  way0_dirty_68 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  way0_dirty_69 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  way0_dirty_70 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  way0_dirty_71 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  way0_dirty_72 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  way0_dirty_73 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  way0_dirty_74 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  way0_dirty_75 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  way0_dirty_76 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  way0_dirty_77 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  way0_dirty_78 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  way0_dirty_79 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  way0_dirty_80 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  way0_dirty_81 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  way0_dirty_82 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  way0_dirty_83 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  way0_dirty_84 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  way0_dirty_85 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  way0_dirty_86 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  way0_dirty_87 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  way0_dirty_88 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  way0_dirty_89 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  way0_dirty_90 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  way0_dirty_91 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  way0_dirty_92 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  way0_dirty_93 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  way0_dirty_94 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  way0_dirty_95 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  way0_dirty_96 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  way0_dirty_97 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  way0_dirty_98 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  way0_dirty_99 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  way0_dirty_100 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  way0_dirty_101 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  way0_dirty_102 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  way0_dirty_103 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  way0_dirty_104 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  way0_dirty_105 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  way0_dirty_106 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  way0_dirty_107 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  way0_dirty_108 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  way0_dirty_109 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  way0_dirty_110 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  way0_dirty_111 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  way0_dirty_112 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  way0_dirty_113 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  way0_dirty_114 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  way0_dirty_115 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  way0_dirty_116 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  way0_dirty_117 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  way0_dirty_118 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  way0_dirty_119 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  way0_dirty_120 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  way0_dirty_121 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  way0_dirty_122 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  way0_dirty_123 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  way0_dirty_124 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  way0_dirty_125 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  way0_dirty_126 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  way0_dirty_127 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  way1_dirty_0 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  way1_dirty_1 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  way1_dirty_2 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  way1_dirty_3 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  way1_dirty_4 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  way1_dirty_5 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  way1_dirty_6 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  way1_dirty_7 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  way1_dirty_8 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  way1_dirty_9 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  way1_dirty_10 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  way1_dirty_11 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  way1_dirty_12 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  way1_dirty_13 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  way1_dirty_14 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  way1_dirty_15 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  way1_dirty_16 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  way1_dirty_17 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  way1_dirty_18 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  way1_dirty_19 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  way1_dirty_20 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  way1_dirty_21 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  way1_dirty_22 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  way1_dirty_23 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  way1_dirty_24 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  way1_dirty_25 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  way1_dirty_26 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  way1_dirty_27 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  way1_dirty_28 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  way1_dirty_29 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  way1_dirty_30 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  way1_dirty_31 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  way1_dirty_32 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  way1_dirty_33 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  way1_dirty_34 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  way1_dirty_35 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  way1_dirty_36 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  way1_dirty_37 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  way1_dirty_38 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  way1_dirty_39 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  way1_dirty_40 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  way1_dirty_41 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  way1_dirty_42 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  way1_dirty_43 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  way1_dirty_44 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  way1_dirty_45 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  way1_dirty_46 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  way1_dirty_47 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  way1_dirty_48 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  way1_dirty_49 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  way1_dirty_50 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  way1_dirty_51 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  way1_dirty_52 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  way1_dirty_53 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  way1_dirty_54 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  way1_dirty_55 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  way1_dirty_56 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  way1_dirty_57 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  way1_dirty_58 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  way1_dirty_59 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  way1_dirty_60 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  way1_dirty_61 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  way1_dirty_62 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  way1_dirty_63 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  way1_dirty_64 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  way1_dirty_65 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  way1_dirty_66 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  way1_dirty_67 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  way1_dirty_68 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  way1_dirty_69 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  way1_dirty_70 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  way1_dirty_71 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  way1_dirty_72 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  way1_dirty_73 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  way1_dirty_74 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  way1_dirty_75 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  way1_dirty_76 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  way1_dirty_77 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  way1_dirty_78 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  way1_dirty_79 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  way1_dirty_80 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  way1_dirty_81 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  way1_dirty_82 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  way1_dirty_83 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  way1_dirty_84 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  way1_dirty_85 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  way1_dirty_86 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  way1_dirty_87 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  way1_dirty_88 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  way1_dirty_89 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  way1_dirty_90 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  way1_dirty_91 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  way1_dirty_92 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  way1_dirty_93 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  way1_dirty_94 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  way1_dirty_95 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  way1_dirty_96 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  way1_dirty_97 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  way1_dirty_98 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  way1_dirty_99 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  way1_dirty_100 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  way1_dirty_101 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  way1_dirty_102 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  way1_dirty_103 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  way1_dirty_104 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  way1_dirty_105 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  way1_dirty_106 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  way1_dirty_107 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  way1_dirty_108 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  way1_dirty_109 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  way1_dirty_110 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  way1_dirty_111 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  way1_dirty_112 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  way1_dirty_113 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  way1_dirty_114 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  way1_dirty_115 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  way1_dirty_116 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  way1_dirty_117 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  way1_dirty_118 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  way1_dirty_119 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  way1_dirty_120 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  way1_dirty_121 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  way1_dirty_122 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  way1_dirty_123 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  way1_dirty_124 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  way1_dirty_125 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  way1_dirty_126 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  way1_dirty_127 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  stage1_sram_addr_reg = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  stage1_sram_cache_reg = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  stage1_sram_wdata_reg = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  stage1_sram_size_reg = _RAND_391[1:0];
  _RAND_392 = {1{`RANDOM}};
  stage1_sram_wr_reg = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  stage1_sram_req_reg = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  stage1_sram_hit0_reg = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  stage1_sram_hit1_reg = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  stage1_sram_valid0_reg = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  stage1_sram_valid1_reg = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  stage1_wstrb_reg = _RAND_398[3:0];
  _RAND_399 = {1{`RANDOM}};
  stage1_sram_phy_addr_reg = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  stage1_exception = _RAND_400[2:0];
  _RAND_401 = {1{`RANDOM}};
  stage2_sram_write_reg = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  stage1_stall_reg = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  write_access_complete_reg = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  stage2_sram_addr_reg = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  stage2_hit0_reg = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  sram_rdata_reg = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  stage2_stall_reg = _RAND_407[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    work_state = 5'h18;
  end
  if (reset) begin
    write_counter = 3'h0;
  end
  if (reset) begin
    read_counter = 3'h0;
  end
  if (reset) begin
    wait_data = 32'h0;
  end
  if (reset) begin
    lru_0 = 1'h0;
  end
  if (reset) begin
    lru_1 = 1'h0;
  end
  if (reset) begin
    lru_2 = 1'h0;
  end
  if (reset) begin
    lru_3 = 1'h0;
  end
  if (reset) begin
    lru_4 = 1'h0;
  end
  if (reset) begin
    lru_5 = 1'h0;
  end
  if (reset) begin
    lru_6 = 1'h0;
  end
  if (reset) begin
    lru_7 = 1'h0;
  end
  if (reset) begin
    lru_8 = 1'h0;
  end
  if (reset) begin
    lru_9 = 1'h0;
  end
  if (reset) begin
    lru_10 = 1'h0;
  end
  if (reset) begin
    lru_11 = 1'h0;
  end
  if (reset) begin
    lru_12 = 1'h0;
  end
  if (reset) begin
    lru_13 = 1'h0;
  end
  if (reset) begin
    lru_14 = 1'h0;
  end
  if (reset) begin
    lru_15 = 1'h0;
  end
  if (reset) begin
    lru_16 = 1'h0;
  end
  if (reset) begin
    lru_17 = 1'h0;
  end
  if (reset) begin
    lru_18 = 1'h0;
  end
  if (reset) begin
    lru_19 = 1'h0;
  end
  if (reset) begin
    lru_20 = 1'h0;
  end
  if (reset) begin
    lru_21 = 1'h0;
  end
  if (reset) begin
    lru_22 = 1'h0;
  end
  if (reset) begin
    lru_23 = 1'h0;
  end
  if (reset) begin
    lru_24 = 1'h0;
  end
  if (reset) begin
    lru_25 = 1'h0;
  end
  if (reset) begin
    lru_26 = 1'h0;
  end
  if (reset) begin
    lru_27 = 1'h0;
  end
  if (reset) begin
    lru_28 = 1'h0;
  end
  if (reset) begin
    lru_29 = 1'h0;
  end
  if (reset) begin
    lru_30 = 1'h0;
  end
  if (reset) begin
    lru_31 = 1'h0;
  end
  if (reset) begin
    lru_32 = 1'h0;
  end
  if (reset) begin
    lru_33 = 1'h0;
  end
  if (reset) begin
    lru_34 = 1'h0;
  end
  if (reset) begin
    lru_35 = 1'h0;
  end
  if (reset) begin
    lru_36 = 1'h0;
  end
  if (reset) begin
    lru_37 = 1'h0;
  end
  if (reset) begin
    lru_38 = 1'h0;
  end
  if (reset) begin
    lru_39 = 1'h0;
  end
  if (reset) begin
    lru_40 = 1'h0;
  end
  if (reset) begin
    lru_41 = 1'h0;
  end
  if (reset) begin
    lru_42 = 1'h0;
  end
  if (reset) begin
    lru_43 = 1'h0;
  end
  if (reset) begin
    lru_44 = 1'h0;
  end
  if (reset) begin
    lru_45 = 1'h0;
  end
  if (reset) begin
    lru_46 = 1'h0;
  end
  if (reset) begin
    lru_47 = 1'h0;
  end
  if (reset) begin
    lru_48 = 1'h0;
  end
  if (reset) begin
    lru_49 = 1'h0;
  end
  if (reset) begin
    lru_50 = 1'h0;
  end
  if (reset) begin
    lru_51 = 1'h0;
  end
  if (reset) begin
    lru_52 = 1'h0;
  end
  if (reset) begin
    lru_53 = 1'h0;
  end
  if (reset) begin
    lru_54 = 1'h0;
  end
  if (reset) begin
    lru_55 = 1'h0;
  end
  if (reset) begin
    lru_56 = 1'h0;
  end
  if (reset) begin
    lru_57 = 1'h0;
  end
  if (reset) begin
    lru_58 = 1'h0;
  end
  if (reset) begin
    lru_59 = 1'h0;
  end
  if (reset) begin
    lru_60 = 1'h0;
  end
  if (reset) begin
    lru_61 = 1'h0;
  end
  if (reset) begin
    lru_62 = 1'h0;
  end
  if (reset) begin
    lru_63 = 1'h0;
  end
  if (reset) begin
    lru_64 = 1'h0;
  end
  if (reset) begin
    lru_65 = 1'h0;
  end
  if (reset) begin
    lru_66 = 1'h0;
  end
  if (reset) begin
    lru_67 = 1'h0;
  end
  if (reset) begin
    lru_68 = 1'h0;
  end
  if (reset) begin
    lru_69 = 1'h0;
  end
  if (reset) begin
    lru_70 = 1'h0;
  end
  if (reset) begin
    lru_71 = 1'h0;
  end
  if (reset) begin
    lru_72 = 1'h0;
  end
  if (reset) begin
    lru_73 = 1'h0;
  end
  if (reset) begin
    lru_74 = 1'h0;
  end
  if (reset) begin
    lru_75 = 1'h0;
  end
  if (reset) begin
    lru_76 = 1'h0;
  end
  if (reset) begin
    lru_77 = 1'h0;
  end
  if (reset) begin
    lru_78 = 1'h0;
  end
  if (reset) begin
    lru_79 = 1'h0;
  end
  if (reset) begin
    lru_80 = 1'h0;
  end
  if (reset) begin
    lru_81 = 1'h0;
  end
  if (reset) begin
    lru_82 = 1'h0;
  end
  if (reset) begin
    lru_83 = 1'h0;
  end
  if (reset) begin
    lru_84 = 1'h0;
  end
  if (reset) begin
    lru_85 = 1'h0;
  end
  if (reset) begin
    lru_86 = 1'h0;
  end
  if (reset) begin
    lru_87 = 1'h0;
  end
  if (reset) begin
    lru_88 = 1'h0;
  end
  if (reset) begin
    lru_89 = 1'h0;
  end
  if (reset) begin
    lru_90 = 1'h0;
  end
  if (reset) begin
    lru_91 = 1'h0;
  end
  if (reset) begin
    lru_92 = 1'h0;
  end
  if (reset) begin
    lru_93 = 1'h0;
  end
  if (reset) begin
    lru_94 = 1'h0;
  end
  if (reset) begin
    lru_95 = 1'h0;
  end
  if (reset) begin
    lru_96 = 1'h0;
  end
  if (reset) begin
    lru_97 = 1'h0;
  end
  if (reset) begin
    lru_98 = 1'h0;
  end
  if (reset) begin
    lru_99 = 1'h0;
  end
  if (reset) begin
    lru_100 = 1'h0;
  end
  if (reset) begin
    lru_101 = 1'h0;
  end
  if (reset) begin
    lru_102 = 1'h0;
  end
  if (reset) begin
    lru_103 = 1'h0;
  end
  if (reset) begin
    lru_104 = 1'h0;
  end
  if (reset) begin
    lru_105 = 1'h0;
  end
  if (reset) begin
    lru_106 = 1'h0;
  end
  if (reset) begin
    lru_107 = 1'h0;
  end
  if (reset) begin
    lru_108 = 1'h0;
  end
  if (reset) begin
    lru_109 = 1'h0;
  end
  if (reset) begin
    lru_110 = 1'h0;
  end
  if (reset) begin
    lru_111 = 1'h0;
  end
  if (reset) begin
    lru_112 = 1'h0;
  end
  if (reset) begin
    lru_113 = 1'h0;
  end
  if (reset) begin
    lru_114 = 1'h0;
  end
  if (reset) begin
    lru_115 = 1'h0;
  end
  if (reset) begin
    lru_116 = 1'h0;
  end
  if (reset) begin
    lru_117 = 1'h0;
  end
  if (reset) begin
    lru_118 = 1'h0;
  end
  if (reset) begin
    lru_119 = 1'h0;
  end
  if (reset) begin
    lru_120 = 1'h0;
  end
  if (reset) begin
    lru_121 = 1'h0;
  end
  if (reset) begin
    lru_122 = 1'h0;
  end
  if (reset) begin
    lru_123 = 1'h0;
  end
  if (reset) begin
    lru_124 = 1'h0;
  end
  if (reset) begin
    lru_125 = 1'h0;
  end
  if (reset) begin
    lru_126 = 1'h0;
  end
  if (reset) begin
    lru_127 = 1'h0;
  end
  if (reset) begin
    way0_dirty_0 = 1'h0;
  end
  if (reset) begin
    way0_dirty_1 = 1'h0;
  end
  if (reset) begin
    way0_dirty_2 = 1'h0;
  end
  if (reset) begin
    way0_dirty_3 = 1'h0;
  end
  if (reset) begin
    way0_dirty_4 = 1'h0;
  end
  if (reset) begin
    way0_dirty_5 = 1'h0;
  end
  if (reset) begin
    way0_dirty_6 = 1'h0;
  end
  if (reset) begin
    way0_dirty_7 = 1'h0;
  end
  if (reset) begin
    way0_dirty_8 = 1'h0;
  end
  if (reset) begin
    way0_dirty_9 = 1'h0;
  end
  if (reset) begin
    way0_dirty_10 = 1'h0;
  end
  if (reset) begin
    way0_dirty_11 = 1'h0;
  end
  if (reset) begin
    way0_dirty_12 = 1'h0;
  end
  if (reset) begin
    way0_dirty_13 = 1'h0;
  end
  if (reset) begin
    way0_dirty_14 = 1'h0;
  end
  if (reset) begin
    way0_dirty_15 = 1'h0;
  end
  if (reset) begin
    way0_dirty_16 = 1'h0;
  end
  if (reset) begin
    way0_dirty_17 = 1'h0;
  end
  if (reset) begin
    way0_dirty_18 = 1'h0;
  end
  if (reset) begin
    way0_dirty_19 = 1'h0;
  end
  if (reset) begin
    way0_dirty_20 = 1'h0;
  end
  if (reset) begin
    way0_dirty_21 = 1'h0;
  end
  if (reset) begin
    way0_dirty_22 = 1'h0;
  end
  if (reset) begin
    way0_dirty_23 = 1'h0;
  end
  if (reset) begin
    way0_dirty_24 = 1'h0;
  end
  if (reset) begin
    way0_dirty_25 = 1'h0;
  end
  if (reset) begin
    way0_dirty_26 = 1'h0;
  end
  if (reset) begin
    way0_dirty_27 = 1'h0;
  end
  if (reset) begin
    way0_dirty_28 = 1'h0;
  end
  if (reset) begin
    way0_dirty_29 = 1'h0;
  end
  if (reset) begin
    way0_dirty_30 = 1'h0;
  end
  if (reset) begin
    way0_dirty_31 = 1'h0;
  end
  if (reset) begin
    way0_dirty_32 = 1'h0;
  end
  if (reset) begin
    way0_dirty_33 = 1'h0;
  end
  if (reset) begin
    way0_dirty_34 = 1'h0;
  end
  if (reset) begin
    way0_dirty_35 = 1'h0;
  end
  if (reset) begin
    way0_dirty_36 = 1'h0;
  end
  if (reset) begin
    way0_dirty_37 = 1'h0;
  end
  if (reset) begin
    way0_dirty_38 = 1'h0;
  end
  if (reset) begin
    way0_dirty_39 = 1'h0;
  end
  if (reset) begin
    way0_dirty_40 = 1'h0;
  end
  if (reset) begin
    way0_dirty_41 = 1'h0;
  end
  if (reset) begin
    way0_dirty_42 = 1'h0;
  end
  if (reset) begin
    way0_dirty_43 = 1'h0;
  end
  if (reset) begin
    way0_dirty_44 = 1'h0;
  end
  if (reset) begin
    way0_dirty_45 = 1'h0;
  end
  if (reset) begin
    way0_dirty_46 = 1'h0;
  end
  if (reset) begin
    way0_dirty_47 = 1'h0;
  end
  if (reset) begin
    way0_dirty_48 = 1'h0;
  end
  if (reset) begin
    way0_dirty_49 = 1'h0;
  end
  if (reset) begin
    way0_dirty_50 = 1'h0;
  end
  if (reset) begin
    way0_dirty_51 = 1'h0;
  end
  if (reset) begin
    way0_dirty_52 = 1'h0;
  end
  if (reset) begin
    way0_dirty_53 = 1'h0;
  end
  if (reset) begin
    way0_dirty_54 = 1'h0;
  end
  if (reset) begin
    way0_dirty_55 = 1'h0;
  end
  if (reset) begin
    way0_dirty_56 = 1'h0;
  end
  if (reset) begin
    way0_dirty_57 = 1'h0;
  end
  if (reset) begin
    way0_dirty_58 = 1'h0;
  end
  if (reset) begin
    way0_dirty_59 = 1'h0;
  end
  if (reset) begin
    way0_dirty_60 = 1'h0;
  end
  if (reset) begin
    way0_dirty_61 = 1'h0;
  end
  if (reset) begin
    way0_dirty_62 = 1'h0;
  end
  if (reset) begin
    way0_dirty_63 = 1'h0;
  end
  if (reset) begin
    way0_dirty_64 = 1'h0;
  end
  if (reset) begin
    way0_dirty_65 = 1'h0;
  end
  if (reset) begin
    way0_dirty_66 = 1'h0;
  end
  if (reset) begin
    way0_dirty_67 = 1'h0;
  end
  if (reset) begin
    way0_dirty_68 = 1'h0;
  end
  if (reset) begin
    way0_dirty_69 = 1'h0;
  end
  if (reset) begin
    way0_dirty_70 = 1'h0;
  end
  if (reset) begin
    way0_dirty_71 = 1'h0;
  end
  if (reset) begin
    way0_dirty_72 = 1'h0;
  end
  if (reset) begin
    way0_dirty_73 = 1'h0;
  end
  if (reset) begin
    way0_dirty_74 = 1'h0;
  end
  if (reset) begin
    way0_dirty_75 = 1'h0;
  end
  if (reset) begin
    way0_dirty_76 = 1'h0;
  end
  if (reset) begin
    way0_dirty_77 = 1'h0;
  end
  if (reset) begin
    way0_dirty_78 = 1'h0;
  end
  if (reset) begin
    way0_dirty_79 = 1'h0;
  end
  if (reset) begin
    way0_dirty_80 = 1'h0;
  end
  if (reset) begin
    way0_dirty_81 = 1'h0;
  end
  if (reset) begin
    way0_dirty_82 = 1'h0;
  end
  if (reset) begin
    way0_dirty_83 = 1'h0;
  end
  if (reset) begin
    way0_dirty_84 = 1'h0;
  end
  if (reset) begin
    way0_dirty_85 = 1'h0;
  end
  if (reset) begin
    way0_dirty_86 = 1'h0;
  end
  if (reset) begin
    way0_dirty_87 = 1'h0;
  end
  if (reset) begin
    way0_dirty_88 = 1'h0;
  end
  if (reset) begin
    way0_dirty_89 = 1'h0;
  end
  if (reset) begin
    way0_dirty_90 = 1'h0;
  end
  if (reset) begin
    way0_dirty_91 = 1'h0;
  end
  if (reset) begin
    way0_dirty_92 = 1'h0;
  end
  if (reset) begin
    way0_dirty_93 = 1'h0;
  end
  if (reset) begin
    way0_dirty_94 = 1'h0;
  end
  if (reset) begin
    way0_dirty_95 = 1'h0;
  end
  if (reset) begin
    way0_dirty_96 = 1'h0;
  end
  if (reset) begin
    way0_dirty_97 = 1'h0;
  end
  if (reset) begin
    way0_dirty_98 = 1'h0;
  end
  if (reset) begin
    way0_dirty_99 = 1'h0;
  end
  if (reset) begin
    way0_dirty_100 = 1'h0;
  end
  if (reset) begin
    way0_dirty_101 = 1'h0;
  end
  if (reset) begin
    way0_dirty_102 = 1'h0;
  end
  if (reset) begin
    way0_dirty_103 = 1'h0;
  end
  if (reset) begin
    way0_dirty_104 = 1'h0;
  end
  if (reset) begin
    way0_dirty_105 = 1'h0;
  end
  if (reset) begin
    way0_dirty_106 = 1'h0;
  end
  if (reset) begin
    way0_dirty_107 = 1'h0;
  end
  if (reset) begin
    way0_dirty_108 = 1'h0;
  end
  if (reset) begin
    way0_dirty_109 = 1'h0;
  end
  if (reset) begin
    way0_dirty_110 = 1'h0;
  end
  if (reset) begin
    way0_dirty_111 = 1'h0;
  end
  if (reset) begin
    way0_dirty_112 = 1'h0;
  end
  if (reset) begin
    way0_dirty_113 = 1'h0;
  end
  if (reset) begin
    way0_dirty_114 = 1'h0;
  end
  if (reset) begin
    way0_dirty_115 = 1'h0;
  end
  if (reset) begin
    way0_dirty_116 = 1'h0;
  end
  if (reset) begin
    way0_dirty_117 = 1'h0;
  end
  if (reset) begin
    way0_dirty_118 = 1'h0;
  end
  if (reset) begin
    way0_dirty_119 = 1'h0;
  end
  if (reset) begin
    way0_dirty_120 = 1'h0;
  end
  if (reset) begin
    way0_dirty_121 = 1'h0;
  end
  if (reset) begin
    way0_dirty_122 = 1'h0;
  end
  if (reset) begin
    way0_dirty_123 = 1'h0;
  end
  if (reset) begin
    way0_dirty_124 = 1'h0;
  end
  if (reset) begin
    way0_dirty_125 = 1'h0;
  end
  if (reset) begin
    way0_dirty_126 = 1'h0;
  end
  if (reset) begin
    way0_dirty_127 = 1'h0;
  end
  if (reset) begin
    way1_dirty_0 = 1'h0;
  end
  if (reset) begin
    way1_dirty_1 = 1'h0;
  end
  if (reset) begin
    way1_dirty_2 = 1'h0;
  end
  if (reset) begin
    way1_dirty_3 = 1'h0;
  end
  if (reset) begin
    way1_dirty_4 = 1'h0;
  end
  if (reset) begin
    way1_dirty_5 = 1'h0;
  end
  if (reset) begin
    way1_dirty_6 = 1'h0;
  end
  if (reset) begin
    way1_dirty_7 = 1'h0;
  end
  if (reset) begin
    way1_dirty_8 = 1'h0;
  end
  if (reset) begin
    way1_dirty_9 = 1'h0;
  end
  if (reset) begin
    way1_dirty_10 = 1'h0;
  end
  if (reset) begin
    way1_dirty_11 = 1'h0;
  end
  if (reset) begin
    way1_dirty_12 = 1'h0;
  end
  if (reset) begin
    way1_dirty_13 = 1'h0;
  end
  if (reset) begin
    way1_dirty_14 = 1'h0;
  end
  if (reset) begin
    way1_dirty_15 = 1'h0;
  end
  if (reset) begin
    way1_dirty_16 = 1'h0;
  end
  if (reset) begin
    way1_dirty_17 = 1'h0;
  end
  if (reset) begin
    way1_dirty_18 = 1'h0;
  end
  if (reset) begin
    way1_dirty_19 = 1'h0;
  end
  if (reset) begin
    way1_dirty_20 = 1'h0;
  end
  if (reset) begin
    way1_dirty_21 = 1'h0;
  end
  if (reset) begin
    way1_dirty_22 = 1'h0;
  end
  if (reset) begin
    way1_dirty_23 = 1'h0;
  end
  if (reset) begin
    way1_dirty_24 = 1'h0;
  end
  if (reset) begin
    way1_dirty_25 = 1'h0;
  end
  if (reset) begin
    way1_dirty_26 = 1'h0;
  end
  if (reset) begin
    way1_dirty_27 = 1'h0;
  end
  if (reset) begin
    way1_dirty_28 = 1'h0;
  end
  if (reset) begin
    way1_dirty_29 = 1'h0;
  end
  if (reset) begin
    way1_dirty_30 = 1'h0;
  end
  if (reset) begin
    way1_dirty_31 = 1'h0;
  end
  if (reset) begin
    way1_dirty_32 = 1'h0;
  end
  if (reset) begin
    way1_dirty_33 = 1'h0;
  end
  if (reset) begin
    way1_dirty_34 = 1'h0;
  end
  if (reset) begin
    way1_dirty_35 = 1'h0;
  end
  if (reset) begin
    way1_dirty_36 = 1'h0;
  end
  if (reset) begin
    way1_dirty_37 = 1'h0;
  end
  if (reset) begin
    way1_dirty_38 = 1'h0;
  end
  if (reset) begin
    way1_dirty_39 = 1'h0;
  end
  if (reset) begin
    way1_dirty_40 = 1'h0;
  end
  if (reset) begin
    way1_dirty_41 = 1'h0;
  end
  if (reset) begin
    way1_dirty_42 = 1'h0;
  end
  if (reset) begin
    way1_dirty_43 = 1'h0;
  end
  if (reset) begin
    way1_dirty_44 = 1'h0;
  end
  if (reset) begin
    way1_dirty_45 = 1'h0;
  end
  if (reset) begin
    way1_dirty_46 = 1'h0;
  end
  if (reset) begin
    way1_dirty_47 = 1'h0;
  end
  if (reset) begin
    way1_dirty_48 = 1'h0;
  end
  if (reset) begin
    way1_dirty_49 = 1'h0;
  end
  if (reset) begin
    way1_dirty_50 = 1'h0;
  end
  if (reset) begin
    way1_dirty_51 = 1'h0;
  end
  if (reset) begin
    way1_dirty_52 = 1'h0;
  end
  if (reset) begin
    way1_dirty_53 = 1'h0;
  end
  if (reset) begin
    way1_dirty_54 = 1'h0;
  end
  if (reset) begin
    way1_dirty_55 = 1'h0;
  end
  if (reset) begin
    way1_dirty_56 = 1'h0;
  end
  if (reset) begin
    way1_dirty_57 = 1'h0;
  end
  if (reset) begin
    way1_dirty_58 = 1'h0;
  end
  if (reset) begin
    way1_dirty_59 = 1'h0;
  end
  if (reset) begin
    way1_dirty_60 = 1'h0;
  end
  if (reset) begin
    way1_dirty_61 = 1'h0;
  end
  if (reset) begin
    way1_dirty_62 = 1'h0;
  end
  if (reset) begin
    way1_dirty_63 = 1'h0;
  end
  if (reset) begin
    way1_dirty_64 = 1'h0;
  end
  if (reset) begin
    way1_dirty_65 = 1'h0;
  end
  if (reset) begin
    way1_dirty_66 = 1'h0;
  end
  if (reset) begin
    way1_dirty_67 = 1'h0;
  end
  if (reset) begin
    way1_dirty_68 = 1'h0;
  end
  if (reset) begin
    way1_dirty_69 = 1'h0;
  end
  if (reset) begin
    way1_dirty_70 = 1'h0;
  end
  if (reset) begin
    way1_dirty_71 = 1'h0;
  end
  if (reset) begin
    way1_dirty_72 = 1'h0;
  end
  if (reset) begin
    way1_dirty_73 = 1'h0;
  end
  if (reset) begin
    way1_dirty_74 = 1'h0;
  end
  if (reset) begin
    way1_dirty_75 = 1'h0;
  end
  if (reset) begin
    way1_dirty_76 = 1'h0;
  end
  if (reset) begin
    way1_dirty_77 = 1'h0;
  end
  if (reset) begin
    way1_dirty_78 = 1'h0;
  end
  if (reset) begin
    way1_dirty_79 = 1'h0;
  end
  if (reset) begin
    way1_dirty_80 = 1'h0;
  end
  if (reset) begin
    way1_dirty_81 = 1'h0;
  end
  if (reset) begin
    way1_dirty_82 = 1'h0;
  end
  if (reset) begin
    way1_dirty_83 = 1'h0;
  end
  if (reset) begin
    way1_dirty_84 = 1'h0;
  end
  if (reset) begin
    way1_dirty_85 = 1'h0;
  end
  if (reset) begin
    way1_dirty_86 = 1'h0;
  end
  if (reset) begin
    way1_dirty_87 = 1'h0;
  end
  if (reset) begin
    way1_dirty_88 = 1'h0;
  end
  if (reset) begin
    way1_dirty_89 = 1'h0;
  end
  if (reset) begin
    way1_dirty_90 = 1'h0;
  end
  if (reset) begin
    way1_dirty_91 = 1'h0;
  end
  if (reset) begin
    way1_dirty_92 = 1'h0;
  end
  if (reset) begin
    way1_dirty_93 = 1'h0;
  end
  if (reset) begin
    way1_dirty_94 = 1'h0;
  end
  if (reset) begin
    way1_dirty_95 = 1'h0;
  end
  if (reset) begin
    way1_dirty_96 = 1'h0;
  end
  if (reset) begin
    way1_dirty_97 = 1'h0;
  end
  if (reset) begin
    way1_dirty_98 = 1'h0;
  end
  if (reset) begin
    way1_dirty_99 = 1'h0;
  end
  if (reset) begin
    way1_dirty_100 = 1'h0;
  end
  if (reset) begin
    way1_dirty_101 = 1'h0;
  end
  if (reset) begin
    way1_dirty_102 = 1'h0;
  end
  if (reset) begin
    way1_dirty_103 = 1'h0;
  end
  if (reset) begin
    way1_dirty_104 = 1'h0;
  end
  if (reset) begin
    way1_dirty_105 = 1'h0;
  end
  if (reset) begin
    way1_dirty_106 = 1'h0;
  end
  if (reset) begin
    way1_dirty_107 = 1'h0;
  end
  if (reset) begin
    way1_dirty_108 = 1'h0;
  end
  if (reset) begin
    way1_dirty_109 = 1'h0;
  end
  if (reset) begin
    way1_dirty_110 = 1'h0;
  end
  if (reset) begin
    way1_dirty_111 = 1'h0;
  end
  if (reset) begin
    way1_dirty_112 = 1'h0;
  end
  if (reset) begin
    way1_dirty_113 = 1'h0;
  end
  if (reset) begin
    way1_dirty_114 = 1'h0;
  end
  if (reset) begin
    way1_dirty_115 = 1'h0;
  end
  if (reset) begin
    way1_dirty_116 = 1'h0;
  end
  if (reset) begin
    way1_dirty_117 = 1'h0;
  end
  if (reset) begin
    way1_dirty_118 = 1'h0;
  end
  if (reset) begin
    way1_dirty_119 = 1'h0;
  end
  if (reset) begin
    way1_dirty_120 = 1'h0;
  end
  if (reset) begin
    way1_dirty_121 = 1'h0;
  end
  if (reset) begin
    way1_dirty_122 = 1'h0;
  end
  if (reset) begin
    way1_dirty_123 = 1'h0;
  end
  if (reset) begin
    way1_dirty_124 = 1'h0;
  end
  if (reset) begin
    way1_dirty_125 = 1'h0;
  end
  if (reset) begin
    way1_dirty_126 = 1'h0;
  end
  if (reset) begin
    way1_dirty_127 = 1'h0;
  end
  if (reset) begin
    stage1_sram_addr_reg = 32'h0;
  end
  if (reset) begin
    stage1_sram_cache_reg = 1'h0;
  end
  if (reset) begin
    stage1_sram_wdata_reg = 32'h0;
  end
  if (reset) begin
    stage1_sram_size_reg = 2'h0;
  end
  if (reset) begin
    stage1_sram_wr_reg = 1'h0;
  end
  if (reset) begin
    stage1_sram_req_reg = 1'h0;
  end
  if (reset) begin
    stage1_sram_hit0_reg = 1'h0;
  end
  if (reset) begin
    stage1_sram_hit1_reg = 1'h0;
  end
  if (reset) begin
    stage1_sram_valid0_reg = 1'h0;
  end
  if (reset) begin
    stage1_sram_valid1_reg = 1'h0;
  end
  if (reset) begin
    stage1_wstrb_reg = 4'h0;
  end
  if (reset) begin
    stage1_sram_phy_addr_reg = 32'h0;
  end
  if (reset) begin
    stage1_exception = 3'h0;
  end
  if (reset) begin
    stage2_sram_write_reg = 1'h0;
  end
  if (reset) begin
    stage1_stall_reg = 1'h0;
  end
  if (reset) begin
    write_access_complete_reg = 1'h0;
  end
  if (reset) begin
    stage2_sram_addr_reg = 32'h0;
  end
  if (reset) begin
    stage2_hit0_reg = 1'h0;
  end
  if (reset) begin
    sram_rdata_reg = 32'h0;
  end
  if (reset) begin
    stage2_stall_reg = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module tlb(
  input         clock,
  input         reset,
  input  [31:0] io_vaddr,
  output [31:0] io_paddr,
  input  [7:0]  io_cp0_asid,
  input  [3:0]  io_tlb_write_index,
  input  [3:0]  io_tlb_read_index,
  input         io_tlb_write_en,
  output [3:0]  io_tlb_search_index,
  output        io_tlb_search_hit,
  output        io_tlb_search_ineffective,
  output        io_tlb_search_has_changed,
  input  [18:0] io_tlb_write_port_vaddr,
  input  [7:0]  io_tlb_write_port_asid,
  input         io_tlb_write_port_g,
  input  [19:0] io_tlb_write_port_paddr_0,
  input  [19:0] io_tlb_write_port_paddr_1,
  input  [2:0]  io_tlb_write_port_c_0,
  input  [2:0]  io_tlb_write_port_c_1,
  input         io_tlb_write_port_d_0,
  input         io_tlb_write_port_d_1,
  input         io_tlb_write_port_v_0,
  input         io_tlb_write_port_v_1,
  output [18:0] io_tlb_read_port_vaddr,
  output [7:0]  io_tlb_read_port_asid,
  output        io_tlb_read_port_g,
  output [19:0] io_tlb_read_port_paddr_0,
  output [19:0] io_tlb_read_port_paddr_1,
  output [2:0]  io_tlb_read_port_c_0,
  output [2:0]  io_tlb_read_port_c_1,
  output        io_tlb_read_port_d_0,
  output        io_tlb_read_port_d_1,
  output        io_tlb_read_port_v_0,
  output        io_tlb_read_port_v_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [95:0] _RAND_2;
  reg [95:0] _RAND_3;
  reg [95:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [95:0] _RAND_6;
  reg [95:0] _RAND_7;
  reg [95:0] _RAND_8;
  reg [95:0] _RAND_9;
  reg [95:0] _RAND_10;
  reg [95:0] _RAND_11;
  reg [95:0] _RAND_12;
  reg [95:0] _RAND_13;
  reg [95:0] _RAND_14;
  reg [95:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [77:0] tlb_reg_0; // @[tlb.scala 85:26]
  reg [77:0] tlb_reg_1; // @[tlb.scala 85:26]
  reg [77:0] tlb_reg_2; // @[tlb.scala 85:26]
  reg [77:0] tlb_reg_3; // @[tlb.scala 85:26]
  reg [77:0] tlb_reg_4; // @[tlb.scala 85:26]
  reg [77:0] tlb_reg_5; // @[tlb.scala 85:26]
  reg [77:0] tlb_reg_6; // @[tlb.scala 85:26]
  reg [77:0] tlb_reg_7; // @[tlb.scala 85:26]
  reg [77:0] tlb_reg_8; // @[tlb.scala 85:26]
  reg [77:0] tlb_reg_9; // @[tlb.scala 85:26]
  reg [77:0] tlb_reg_10; // @[tlb.scala 85:26]
  reg [77:0] tlb_reg_11; // @[tlb.scala 85:26]
  reg [77:0] tlb_reg_12; // @[tlb.scala 85:26]
  reg [77:0] tlb_reg_13; // @[tlb.scala 85:26]
  reg [77:0] tlb_reg_14; // @[tlb.scala 85:26]
  reg [77:0] tlb_reg_15; // @[tlb.scala 85:26]
  wire  tlb_search_answer_0 = tlb_reg_0[77:59] == io_vaddr[31:13]; // @[tlb.scala 90:54]
  wire  tlb_search_answer_1 = tlb_reg_1[77:59] == io_vaddr[31:13]; // @[tlb.scala 90:54]
  wire  tlb_search_answer_2 = tlb_reg_2[77:59] == io_vaddr[31:13]; // @[tlb.scala 90:54]
  wire  tlb_search_answer_3 = tlb_reg_3[77:59] == io_vaddr[31:13]; // @[tlb.scala 90:54]
  wire  tlb_search_answer_4 = tlb_reg_4[77:59] == io_vaddr[31:13]; // @[tlb.scala 90:54]
  wire  tlb_search_answer_5 = tlb_reg_5[77:59] == io_vaddr[31:13]; // @[tlb.scala 90:54]
  wire  tlb_search_answer_6 = tlb_reg_6[77:59] == io_vaddr[31:13]; // @[tlb.scala 90:54]
  wire  tlb_search_answer_7 = tlb_reg_7[77:59] == io_vaddr[31:13]; // @[tlb.scala 90:54]
  wire  tlb_search_answer_8 = tlb_reg_8[77:59] == io_vaddr[31:13]; // @[tlb.scala 90:54]
  wire  tlb_search_answer_9 = tlb_reg_9[77:59] == io_vaddr[31:13]; // @[tlb.scala 90:54]
  wire  tlb_search_answer_10 = tlb_reg_10[77:59] == io_vaddr[31:13]; // @[tlb.scala 90:54]
  wire  tlb_search_answer_11 = tlb_reg_11[77:59] == io_vaddr[31:13]; // @[tlb.scala 90:54]
  wire  tlb_search_answer_12 = tlb_reg_12[77:59] == io_vaddr[31:13]; // @[tlb.scala 90:54]
  wire  tlb_search_answer_13 = tlb_reg_13[77:59] == io_vaddr[31:13]; // @[tlb.scala 90:54]
  wire  tlb_search_answer_14 = tlb_reg_14[77:59] == io_vaddr[31:13]; // @[tlb.scala 90:54]
  wire  tlb_search_answer_15 = tlb_reg_15[77:59] == io_vaddr[31:13]; // @[tlb.scala 90:54]
  wire [77:0] _tlb_search_value_T = tlb_search_answer_0 ? tlb_reg_0 : 78'h0; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_1 = tlb_search_answer_1 ? tlb_reg_1 : 78'h0; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_2 = tlb_search_answer_2 ? tlb_reg_2 : 78'h0; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_3 = tlb_search_answer_3 ? tlb_reg_3 : 78'h0; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_4 = tlb_search_answer_4 ? tlb_reg_4 : 78'h0; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_5 = tlb_search_answer_5 ? tlb_reg_5 : 78'h0; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_6 = tlb_search_answer_6 ? tlb_reg_6 : 78'h0; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_7 = tlb_search_answer_7 ? tlb_reg_7 : 78'h0; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_8 = tlb_search_answer_8 ? tlb_reg_8 : 78'h0; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_9 = tlb_search_answer_9 ? tlb_reg_9 : 78'h0; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_10 = tlb_search_answer_10 ? tlb_reg_10 : 78'h0; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_11 = tlb_search_answer_11 ? tlb_reg_11 : 78'h0; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_12 = tlb_search_answer_12 ? tlb_reg_12 : 78'h0; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_13 = tlb_search_answer_13 ? tlb_reg_13 : 78'h0; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_14 = tlb_search_answer_14 ? tlb_reg_14 : 78'h0; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_15 = tlb_search_answer_15 ? tlb_reg_15 : 78'h0; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_16 = _tlb_search_value_T | _tlb_search_value_T_1; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_17 = _tlb_search_value_T_16 | _tlb_search_value_T_2; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_18 = _tlb_search_value_T_17 | _tlb_search_value_T_3; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_19 = _tlb_search_value_T_18 | _tlb_search_value_T_4; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_20 = _tlb_search_value_T_19 | _tlb_search_value_T_5; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_21 = _tlb_search_value_T_20 | _tlb_search_value_T_6; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_22 = _tlb_search_value_T_21 | _tlb_search_value_T_7; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_23 = _tlb_search_value_T_22 | _tlb_search_value_T_8; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_24 = _tlb_search_value_T_23 | _tlb_search_value_T_9; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_25 = _tlb_search_value_T_24 | _tlb_search_value_T_10; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_26 = _tlb_search_value_T_25 | _tlb_search_value_T_11; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_27 = _tlb_search_value_T_26 | _tlb_search_value_T_12; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_28 = _tlb_search_value_T_27 | _tlb_search_value_T_13; // @[Mux.scala 27:73]
  wire [77:0] _tlb_search_value_T_29 = _tlb_search_value_T_28 | _tlb_search_value_T_14; // @[Mux.scala 27:73]
  wire [77:0] tlb_search_value = _tlb_search_value_T_29 | _tlb_search_value_T_15; // @[Mux.scala 27:73]
  wire [7:0] tlb_search_hit_lo = {tlb_search_answer_7,tlb_search_answer_6,tlb_search_answer_5,tlb_search_answer_4,
    tlb_search_answer_3,tlb_search_answer_2,tlb_search_answer_1,tlb_search_answer_0}; // @[tlb.scala 102:41]
  wire [15:0] _tlb_search_hit_T = {tlb_search_answer_15,tlb_search_answer_14,tlb_search_answer_13,tlb_search_answer_12,
    tlb_search_answer_11,tlb_search_answer_10,tlb_search_answer_9,tlb_search_answer_8,tlb_search_hit_lo}; // @[tlb.scala 102:41]
  wire  tlb_search_hit = _tlb_search_hit_T != 16'h0 & (tlb_search_value[58:51] == io_cp0_asid | tlb_search_value[50]); // @[tlb.scala 102:56]
  wire [19:0] tlb_search_phy = io_vaddr[12] ? tlb_search_value[24:5] : tlb_search_value[49:30]; // @[tlb.scala 105:26]
  wire [25:0] tlb_reg_lo = {io_tlb_write_port_v_0,io_tlb_write_port_paddr_1,io_tlb_write_port_c_1,io_tlb_write_port_d_1,
    io_tlb_write_port_v_1}; // @[Cat.scala 31:58]
  wire [77:0] _tlb_reg_T = {io_tlb_write_port_vaddr,io_tlb_write_port_asid,io_tlb_write_port_g,io_tlb_write_port_paddr_0
    ,io_tlb_write_port_c_0,io_tlb_write_port_d_0,tlb_reg_lo}; // @[Cat.scala 31:58]
  wire [77:0] _GEN_1 = 4'h1 == io_tlb_write_index ? tlb_reg_1 : tlb_reg_0; // @[tlb.scala 107:{39,39}]
  wire [77:0] _GEN_2 = 4'h2 == io_tlb_write_index ? tlb_reg_2 : _GEN_1; // @[tlb.scala 107:{39,39}]
  wire [77:0] _GEN_3 = 4'h3 == io_tlb_write_index ? tlb_reg_3 : _GEN_2; // @[tlb.scala 107:{39,39}]
  wire [77:0] _GEN_4 = 4'h4 == io_tlb_write_index ? tlb_reg_4 : _GEN_3; // @[tlb.scala 107:{39,39}]
  wire [77:0] _GEN_5 = 4'h5 == io_tlb_write_index ? tlb_reg_5 : _GEN_4; // @[tlb.scala 107:{39,39}]
  wire [77:0] _GEN_6 = 4'h6 == io_tlb_write_index ? tlb_reg_6 : _GEN_5; // @[tlb.scala 107:{39,39}]
  wire [77:0] _GEN_7 = 4'h7 == io_tlb_write_index ? tlb_reg_7 : _GEN_6; // @[tlb.scala 107:{39,39}]
  wire [77:0] _GEN_8 = 4'h8 == io_tlb_write_index ? tlb_reg_8 : _GEN_7; // @[tlb.scala 107:{39,39}]
  wire [77:0] _GEN_9 = 4'h9 == io_tlb_write_index ? tlb_reg_9 : _GEN_8; // @[tlb.scala 107:{39,39}]
  wire [77:0] _GEN_10 = 4'ha == io_tlb_write_index ? tlb_reg_10 : _GEN_9; // @[tlb.scala 107:{39,39}]
  wire [77:0] _GEN_11 = 4'hb == io_tlb_write_index ? tlb_reg_11 : _GEN_10; // @[tlb.scala 107:{39,39}]
  wire [77:0] _GEN_12 = 4'hc == io_tlb_write_index ? tlb_reg_12 : _GEN_11; // @[tlb.scala 107:{39,39}]
  wire [77:0] _GEN_13 = 4'hd == io_tlb_write_index ? tlb_reg_13 : _GEN_12; // @[tlb.scala 107:{39,39}]
  wire  _io_tlb_search_ineffective_T_5 = io_vaddr[12] ? tlb_search_value[0] : tlb_search_value[25]; // @[tlb.scala 115:58]
  wire  _io_tlb_search_has_changed_T_12 = io_vaddr[12] ? tlb_search_value[1] : tlb_search_value[26]; // @[tlb.scala 117:13]
  wire  _io_tlb_search_has_changed_T_13 = ~_io_tlb_search_has_changed_T_12; // @[tlb.scala 117:9]
  wire [77:0] _GEN_33 = 4'h1 == io_tlb_read_index ? tlb_reg_1 : tlb_reg_0; // @[tlb.scala 61:{47,47}]
  wire [77:0] _GEN_34 = 4'h2 == io_tlb_read_index ? tlb_reg_2 : _GEN_33; // @[tlb.scala 61:{47,47}]
  wire [77:0] _GEN_35 = 4'h3 == io_tlb_read_index ? tlb_reg_3 : _GEN_34; // @[tlb.scala 61:{47,47}]
  wire [77:0] _GEN_36 = 4'h4 == io_tlb_read_index ? tlb_reg_4 : _GEN_35; // @[tlb.scala 61:{47,47}]
  wire [77:0] _GEN_37 = 4'h5 == io_tlb_read_index ? tlb_reg_5 : _GEN_36; // @[tlb.scala 61:{47,47}]
  wire [77:0] _GEN_38 = 4'h6 == io_tlb_read_index ? tlb_reg_6 : _GEN_37; // @[tlb.scala 61:{47,47}]
  wire [77:0] _GEN_39 = 4'h7 == io_tlb_read_index ? tlb_reg_7 : _GEN_38; // @[tlb.scala 61:{47,47}]
  wire [77:0] _GEN_40 = 4'h8 == io_tlb_read_index ? tlb_reg_8 : _GEN_39; // @[tlb.scala 61:{47,47}]
  wire [77:0] _GEN_41 = 4'h9 == io_tlb_read_index ? tlb_reg_9 : _GEN_40; // @[tlb.scala 61:{47,47}]
  wire [77:0] _GEN_42 = 4'ha == io_tlb_read_index ? tlb_reg_10 : _GEN_41; // @[tlb.scala 61:{47,47}]
  wire [77:0] _GEN_43 = 4'hb == io_tlb_read_index ? tlb_reg_11 : _GEN_42; // @[tlb.scala 61:{47,47}]
  wire [77:0] _GEN_44 = 4'hc == io_tlb_read_index ? tlb_reg_12 : _GEN_43; // @[tlb.scala 61:{47,47}]
  wire [77:0] _GEN_45 = 4'hd == io_tlb_read_index ? tlb_reg_13 : _GEN_44; // @[tlb.scala 61:{47,47}]
  wire [77:0] _GEN_46 = 4'he == io_tlb_read_index ? tlb_reg_14 : _GEN_45; // @[tlb.scala 61:{47,47}]
  wire [77:0] _GEN_47 = 4'hf == io_tlb_read_index ? tlb_reg_15 : _GEN_46; // @[tlb.scala 61:{47,47}]
  wire [1:0] _io_tlb_search_index_T_2 = tlb_search_answer_2 ? 2'h2 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_tlb_search_index_T_3 = tlb_search_answer_3 ? 2'h3 : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_tlb_search_index_T_4 = tlb_search_answer_4 ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_tlb_search_index_T_5 = tlb_search_answer_5 ? 3'h5 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_tlb_search_index_T_6 = tlb_search_answer_6 ? 3'h6 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_tlb_search_index_T_7 = tlb_search_answer_7 ? 3'h7 : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_tlb_search_index_T_8 = tlb_search_answer_8 ? 4'h8 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_tlb_search_index_T_9 = tlb_search_answer_9 ? 4'h9 : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_tlb_search_index_T_10 = tlb_search_answer_10 ? 4'ha : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_tlb_search_index_T_11 = tlb_search_answer_11 ? 4'hb : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_tlb_search_index_T_12 = tlb_search_answer_12 ? 4'hc : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_tlb_search_index_T_13 = tlb_search_answer_13 ? 4'hd : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_tlb_search_index_T_14 = tlb_search_answer_14 ? 4'he : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_tlb_search_index_T_15 = tlb_search_answer_15 ? 4'hf : 4'h0; // @[Mux.scala 27:73]
  wire [1:0] _GEN_48 = {{1'd0}, tlb_search_answer_1}; // @[Mux.scala 27:73]
  wire [1:0] _io_tlb_search_index_T_17 = _GEN_48 | _io_tlb_search_index_T_2; // @[Mux.scala 27:73]
  wire [1:0] _io_tlb_search_index_T_18 = _io_tlb_search_index_T_17 | _io_tlb_search_index_T_3; // @[Mux.scala 27:73]
  wire [2:0] _GEN_49 = {{1'd0}, _io_tlb_search_index_T_18}; // @[Mux.scala 27:73]
  wire [2:0] _io_tlb_search_index_T_19 = _GEN_49 | _io_tlb_search_index_T_4; // @[Mux.scala 27:73]
  wire [2:0] _io_tlb_search_index_T_20 = _io_tlb_search_index_T_19 | _io_tlb_search_index_T_5; // @[Mux.scala 27:73]
  wire [2:0] _io_tlb_search_index_T_21 = _io_tlb_search_index_T_20 | _io_tlb_search_index_T_6; // @[Mux.scala 27:73]
  wire [2:0] _io_tlb_search_index_T_22 = _io_tlb_search_index_T_21 | _io_tlb_search_index_T_7; // @[Mux.scala 27:73]
  wire [3:0] _GEN_50 = {{1'd0}, _io_tlb_search_index_T_22}; // @[Mux.scala 27:73]
  wire [3:0] _io_tlb_search_index_T_23 = _GEN_50 | _io_tlb_search_index_T_8; // @[Mux.scala 27:73]
  wire [3:0] _io_tlb_search_index_T_24 = _io_tlb_search_index_T_23 | _io_tlb_search_index_T_9; // @[Mux.scala 27:73]
  wire [3:0] _io_tlb_search_index_T_25 = _io_tlb_search_index_T_24 | _io_tlb_search_index_T_10; // @[Mux.scala 27:73]
  wire [3:0] _io_tlb_search_index_T_26 = _io_tlb_search_index_T_25 | _io_tlb_search_index_T_11; // @[Mux.scala 27:73]
  wire [3:0] _io_tlb_search_index_T_27 = _io_tlb_search_index_T_26 | _io_tlb_search_index_T_12; // @[Mux.scala 27:73]
  wire [3:0] _io_tlb_search_index_T_28 = _io_tlb_search_index_T_27 | _io_tlb_search_index_T_13; // @[Mux.scala 27:73]
  wire [3:0] _io_tlb_search_index_T_29 = _io_tlb_search_index_T_28 | _io_tlb_search_index_T_14; // @[Mux.scala 27:73]
  assign io_paddr = {tlb_search_phy,io_vaddr[11:0]}; // @[Cat.scala 31:58]
  assign io_tlb_search_index = _io_tlb_search_index_T_29 | _io_tlb_search_index_T_15; // @[Mux.scala 27:73]
  assign io_tlb_search_hit = _tlb_search_hit_T != 16'h0 & (tlb_search_value[58:51] == io_cp0_asid | tlb_search_value[50]
    ); // @[tlb.scala 102:56]
  assign io_tlb_search_ineffective = tlb_search_hit & ~_io_tlb_search_ineffective_T_5; // @[tlb.scala 115:50]
  assign io_tlb_search_has_changed = tlb_search_hit & _io_tlb_search_ineffective_T_5 & _io_tlb_search_has_changed_T_13; // @[tlb.scala 116:132]
  assign io_tlb_read_port_vaddr = _GEN_47[77:59]; // @[tlb.scala 67:43]
  assign io_tlb_read_port_asid = _GEN_47[58:51]; // @[tlb.scala 66:43]
  assign io_tlb_read_port_g = _GEN_47[50]; // @[tlb.scala 65:41]
  assign io_tlb_read_port_paddr_0 = _GEN_47[49:30]; // @[tlb.scala 64:47]
  assign io_tlb_read_port_paddr_1 = _GEN_47[24:5]; // @[tlb.scala 62:47]
  assign io_tlb_read_port_c_0 = _GEN_47[29:27]; // @[tlb.scala 125:57]
  assign io_tlb_read_port_c_1 = _GEN_47[4:2]; // @[tlb.scala 122:57]
  assign io_tlb_read_port_d_0 = _GEN_47[26]; // @[tlb.scala 124:57]
  assign io_tlb_read_port_d_1 = _GEN_47[1]; // @[tlb.scala 121:57]
  assign io_tlb_read_port_v_0 = _GEN_47[25]; // @[tlb.scala 123:57]
  assign io_tlb_read_port_v_1 = _GEN_47[0]; // @[tlb.scala 120:57]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[tlb.scala 107:33]
      tlb_reg_0 <= 78'h0; // @[tlb.scala 107:{39,39,39,39,39}]
    end else if (4'h0 == io_tlb_write_index) begin // @[tlb.scala 85:26]
      if (io_tlb_write_en) begin
        tlb_reg_0 <= _tlb_reg_T;
      end else if (4'hf == io_tlb_write_index) begin
        tlb_reg_0 <= tlb_reg_15;
      end else if (4'he == io_tlb_write_index) begin
        tlb_reg_0 <= tlb_reg_14;
      end else begin
        tlb_reg_0 <= _GEN_13;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[tlb.scala 107:33]
      tlb_reg_1 <= 78'h0; // @[tlb.scala 107:{39,39,39,39,39}]
    end else if (4'h1 == io_tlb_write_index) begin // @[tlb.scala 85:26]
      if (io_tlb_write_en) begin
        tlb_reg_1 <= _tlb_reg_T;
      end else if (4'hf == io_tlb_write_index) begin
        tlb_reg_1 <= tlb_reg_15;
      end else if (4'he == io_tlb_write_index) begin
        tlb_reg_1 <= tlb_reg_14;
      end else begin
        tlb_reg_1 <= _GEN_13;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[tlb.scala 107:33]
      tlb_reg_2 <= 78'h0; // @[tlb.scala 107:{39,39,39,39,39}]
    end else if (4'h2 == io_tlb_write_index) begin // @[tlb.scala 85:26]
      if (io_tlb_write_en) begin
        tlb_reg_2 <= _tlb_reg_T;
      end else if (4'hf == io_tlb_write_index) begin
        tlb_reg_2 <= tlb_reg_15;
      end else if (4'he == io_tlb_write_index) begin
        tlb_reg_2 <= tlb_reg_14;
      end else begin
        tlb_reg_2 <= _GEN_13;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[tlb.scala 107:33]
      tlb_reg_3 <= 78'h0; // @[tlb.scala 107:{39,39,39,39,39}]
    end else if (4'h3 == io_tlb_write_index) begin // @[tlb.scala 85:26]
      if (io_tlb_write_en) begin
        tlb_reg_3 <= _tlb_reg_T;
      end else if (4'hf == io_tlb_write_index) begin
        tlb_reg_3 <= tlb_reg_15;
      end else if (4'he == io_tlb_write_index) begin
        tlb_reg_3 <= tlb_reg_14;
      end else begin
        tlb_reg_3 <= _GEN_13;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[tlb.scala 107:33]
      tlb_reg_4 <= 78'h0; // @[tlb.scala 107:{39,39,39,39,39}]
    end else if (4'h4 == io_tlb_write_index) begin // @[tlb.scala 85:26]
      if (io_tlb_write_en) begin
        tlb_reg_4 <= _tlb_reg_T;
      end else if (4'hf == io_tlb_write_index) begin
        tlb_reg_4 <= tlb_reg_15;
      end else if (4'he == io_tlb_write_index) begin
        tlb_reg_4 <= tlb_reg_14;
      end else begin
        tlb_reg_4 <= _GEN_13;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[tlb.scala 107:33]
      tlb_reg_5 <= 78'h0; // @[tlb.scala 107:{39,39,39,39,39}]
    end else if (4'h5 == io_tlb_write_index) begin // @[tlb.scala 85:26]
      if (io_tlb_write_en) begin
        tlb_reg_5 <= _tlb_reg_T;
      end else if (4'hf == io_tlb_write_index) begin
        tlb_reg_5 <= tlb_reg_15;
      end else if (4'he == io_tlb_write_index) begin
        tlb_reg_5 <= tlb_reg_14;
      end else begin
        tlb_reg_5 <= _GEN_13;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[tlb.scala 107:33]
      tlb_reg_6 <= 78'h0; // @[tlb.scala 107:{39,39,39,39,39}]
    end else if (4'h6 == io_tlb_write_index) begin // @[tlb.scala 85:26]
      if (io_tlb_write_en) begin
        tlb_reg_6 <= _tlb_reg_T;
      end else if (4'hf == io_tlb_write_index) begin
        tlb_reg_6 <= tlb_reg_15;
      end else if (4'he == io_tlb_write_index) begin
        tlb_reg_6 <= tlb_reg_14;
      end else begin
        tlb_reg_6 <= _GEN_13;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[tlb.scala 107:33]
      tlb_reg_7 <= 78'h0; // @[tlb.scala 107:{39,39,39,39,39}]
    end else if (4'h7 == io_tlb_write_index) begin // @[tlb.scala 85:26]
      if (io_tlb_write_en) begin
        tlb_reg_7 <= _tlb_reg_T;
      end else if (4'hf == io_tlb_write_index) begin
        tlb_reg_7 <= tlb_reg_15;
      end else if (4'he == io_tlb_write_index) begin
        tlb_reg_7 <= tlb_reg_14;
      end else begin
        tlb_reg_7 <= _GEN_13;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[tlb.scala 107:33]
      tlb_reg_8 <= 78'h0; // @[tlb.scala 107:{39,39,39,39,39}]
    end else if (4'h8 == io_tlb_write_index) begin // @[tlb.scala 85:26]
      if (io_tlb_write_en) begin
        tlb_reg_8 <= _tlb_reg_T;
      end else if (4'hf == io_tlb_write_index) begin
        tlb_reg_8 <= tlb_reg_15;
      end else if (4'he == io_tlb_write_index) begin
        tlb_reg_8 <= tlb_reg_14;
      end else begin
        tlb_reg_8 <= _GEN_13;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[tlb.scala 107:33]
      tlb_reg_9 <= 78'h0; // @[tlb.scala 107:{39,39,39,39,39}]
    end else if (4'h9 == io_tlb_write_index) begin // @[tlb.scala 85:26]
      if (io_tlb_write_en) begin
        tlb_reg_9 <= _tlb_reg_T;
      end else if (4'hf == io_tlb_write_index) begin
        tlb_reg_9 <= tlb_reg_15;
      end else if (4'he == io_tlb_write_index) begin
        tlb_reg_9 <= tlb_reg_14;
      end else begin
        tlb_reg_9 <= _GEN_13;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[tlb.scala 107:33]
      tlb_reg_10 <= 78'h0; // @[tlb.scala 107:{39,39,39,39,39}]
    end else if (4'ha == io_tlb_write_index) begin // @[tlb.scala 85:26]
      if (io_tlb_write_en) begin
        tlb_reg_10 <= _tlb_reg_T;
      end else if (4'hf == io_tlb_write_index) begin
        tlb_reg_10 <= tlb_reg_15;
      end else if (4'he == io_tlb_write_index) begin
        tlb_reg_10 <= tlb_reg_14;
      end else begin
        tlb_reg_10 <= _GEN_13;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[tlb.scala 107:33]
      tlb_reg_11 <= 78'h0; // @[tlb.scala 107:{39,39,39,39,39}]
    end else if (4'hb == io_tlb_write_index) begin // @[tlb.scala 85:26]
      if (io_tlb_write_en) begin
        tlb_reg_11 <= _tlb_reg_T;
      end else if (4'hf == io_tlb_write_index) begin
        tlb_reg_11 <= tlb_reg_15;
      end else if (4'he == io_tlb_write_index) begin
        tlb_reg_11 <= tlb_reg_14;
      end else begin
        tlb_reg_11 <= _GEN_13;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[tlb.scala 107:33]
      tlb_reg_12 <= 78'h0; // @[tlb.scala 107:{39,39,39,39,39}]
    end else if (4'hc == io_tlb_write_index) begin // @[tlb.scala 85:26]
      if (io_tlb_write_en) begin
        tlb_reg_12 <= _tlb_reg_T;
      end else if (4'hf == io_tlb_write_index) begin
        tlb_reg_12 <= tlb_reg_15;
      end else if (4'he == io_tlb_write_index) begin
        tlb_reg_12 <= tlb_reg_14;
      end else begin
        tlb_reg_12 <= _GEN_13;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[tlb.scala 107:33]
      tlb_reg_13 <= 78'h0; // @[tlb.scala 107:{39,39,39,39,39}]
    end else if (4'hd == io_tlb_write_index) begin // @[tlb.scala 85:26]
      if (io_tlb_write_en) begin
        tlb_reg_13 <= _tlb_reg_T;
      end else if (4'hf == io_tlb_write_index) begin
        tlb_reg_13 <= tlb_reg_15;
      end else if (4'he == io_tlb_write_index) begin
        tlb_reg_13 <= tlb_reg_14;
      end else begin
        tlb_reg_13 <= _GEN_13;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[tlb.scala 107:33]
      tlb_reg_14 <= 78'h0; // @[tlb.scala 107:{39,39,39,39,39}]
    end else if (4'he == io_tlb_write_index) begin // @[tlb.scala 85:26]
      if (io_tlb_write_en) begin
        tlb_reg_14 <= _tlb_reg_T;
      end else if (4'hf == io_tlb_write_index) begin
        tlb_reg_14 <= tlb_reg_15;
      end else if (!(4'he == io_tlb_write_index)) begin
        tlb_reg_14 <= _GEN_13;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[tlb.scala 107:33]
      tlb_reg_15 <= 78'h0; // @[tlb.scala 107:{39,39,39,39,39}]
    end else if (4'hf == io_tlb_write_index) begin // @[tlb.scala 85:26]
      if (io_tlb_write_en) begin
        tlb_reg_15 <= _tlb_reg_T;
      end else if (!(4'hf == io_tlb_write_index)) begin
        if (4'he == io_tlb_write_index) begin
          tlb_reg_15 <= tlb_reg_14;
        end else begin
          tlb_reg_15 <= _GEN_13;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  tlb_reg_0 = _RAND_0[77:0];
  _RAND_1 = {3{`RANDOM}};
  tlb_reg_1 = _RAND_1[77:0];
  _RAND_2 = {3{`RANDOM}};
  tlb_reg_2 = _RAND_2[77:0];
  _RAND_3 = {3{`RANDOM}};
  tlb_reg_3 = _RAND_3[77:0];
  _RAND_4 = {3{`RANDOM}};
  tlb_reg_4 = _RAND_4[77:0];
  _RAND_5 = {3{`RANDOM}};
  tlb_reg_5 = _RAND_5[77:0];
  _RAND_6 = {3{`RANDOM}};
  tlb_reg_6 = _RAND_6[77:0];
  _RAND_7 = {3{`RANDOM}};
  tlb_reg_7 = _RAND_7[77:0];
  _RAND_8 = {3{`RANDOM}};
  tlb_reg_8 = _RAND_8[77:0];
  _RAND_9 = {3{`RANDOM}};
  tlb_reg_9 = _RAND_9[77:0];
  _RAND_10 = {3{`RANDOM}};
  tlb_reg_10 = _RAND_10[77:0];
  _RAND_11 = {3{`RANDOM}};
  tlb_reg_11 = _RAND_11[77:0];
  _RAND_12 = {3{`RANDOM}};
  tlb_reg_12 = _RAND_12[77:0];
  _RAND_13 = {3{`RANDOM}};
  tlb_reg_13 = _RAND_13[77:0];
  _RAND_14 = {3{`RANDOM}};
  tlb_reg_14 = _RAND_14[77:0];
  _RAND_15 = {3{`RANDOM}};
  tlb_reg_15 = _RAND_15[77:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    tlb_reg_0 = 78'h0;
  end
  if (reset) begin
    tlb_reg_1 = 78'h0;
  end
  if (reset) begin
    tlb_reg_2 = 78'h0;
  end
  if (reset) begin
    tlb_reg_3 = 78'h0;
  end
  if (reset) begin
    tlb_reg_4 = 78'h0;
  end
  if (reset) begin
    tlb_reg_5 = 78'h0;
  end
  if (reset) begin
    tlb_reg_6 = 78'h0;
  end
  if (reset) begin
    tlb_reg_7 = 78'h0;
  end
  if (reset) begin
    tlb_reg_8 = 78'h0;
  end
  if (reset) begin
    tlb_reg_9 = 78'h0;
  end
  if (reset) begin
    tlb_reg_10 = 78'h0;
  end
  if (reset) begin
    tlb_reg_11 = 78'h0;
  end
  if (reset) begin
    tlb_reg_12 = 78'h0;
  end
  if (reset) begin
    tlb_reg_13 = 78'h0;
  end
  if (reset) begin
    tlb_reg_14 = 78'h0;
  end
  if (reset) begin
    tlb_reg_15 = 78'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module double_ports_tlb_for_inst_and_data(
  input         clock,
  input         reset,
  input  [7:0]  io_cp0_asid,
  input  [3:0]  io_tlb_write_index,
  input  [3:0]  io_tlb_read_index,
  input         io_tlb_write_en,
  output [3:0]  io_tlb_search_index,
  output        io_tlb_search_hit,
  output        io_tlb_dirty_exception,
  input  [18:0] io_tlb_write_port_vaddr,
  input  [7:0]  io_tlb_write_port_asid,
  input         io_tlb_write_port_g,
  input  [19:0] io_tlb_write_port_paddr_0,
  input  [19:0] io_tlb_write_port_paddr_1,
  input  [2:0]  io_tlb_write_port_c_0,
  input  [2:0]  io_tlb_write_port_c_1,
  input         io_tlb_write_port_d_0,
  input         io_tlb_write_port_d_1,
  input         io_tlb_write_port_v_0,
  input         io_tlb_write_port_v_1,
  output [18:0] io_tlb_read_port_vaddr,
  output [7:0]  io_tlb_read_port_asid,
  output        io_tlb_read_port_g,
  output [19:0] io_tlb_read_port_paddr_0,
  output [19:0] io_tlb_read_port_paddr_1,
  output [2:0]  io_tlb_read_port_c_0,
  output [2:0]  io_tlb_read_port_c_1,
  output        io_tlb_read_port_d_0,
  output        io_tlb_read_port_d_1,
  output        io_tlb_read_port_v_0,
  output        io_tlb_read_port_v_1,
  input  [31:0] io_icache_port_vaddr,
  output [31:0] io_icache_port_paddr,
  input         io_icache_port_req,
  output        io_icache_port_tlb_search_not_hit_exception,
  output        io_icache_port_tlb_search_ineffective_exception,
  input  [31:0] io_dcache_port_vaddr,
  output [31:0] io_dcache_port_paddr,
  input         io_dcache_port_req,
  input         io_dcache_port_wr,
  output        io_dcache_port_tlb_search_not_hit_exception,
  output        io_dcache_port_tlb_search_ineffective_exception
);
  wire  tlb_clock; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire  tlb_reset; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [31:0] tlb_io_vaddr; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [31:0] tlb_io_paddr; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [7:0] tlb_io_cp0_asid; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [3:0] tlb_io_tlb_write_index; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [3:0] tlb_io_tlb_read_index; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire  tlb_io_tlb_write_en; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [3:0] tlb_io_tlb_search_index; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire  tlb_io_tlb_search_hit; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire  tlb_io_tlb_search_ineffective; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire  tlb_io_tlb_search_has_changed; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [18:0] tlb_io_tlb_write_port_vaddr; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [7:0] tlb_io_tlb_write_port_asid; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire  tlb_io_tlb_write_port_g; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [19:0] tlb_io_tlb_write_port_paddr_0; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [19:0] tlb_io_tlb_write_port_paddr_1; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [2:0] tlb_io_tlb_write_port_c_0; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [2:0] tlb_io_tlb_write_port_c_1; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire  tlb_io_tlb_write_port_d_0; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire  tlb_io_tlb_write_port_d_1; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire  tlb_io_tlb_write_port_v_0; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire  tlb_io_tlb_write_port_v_1; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [18:0] tlb_io_tlb_read_port_vaddr; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [7:0] tlb_io_tlb_read_port_asid; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire  tlb_io_tlb_read_port_g; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [19:0] tlb_io_tlb_read_port_paddr_0; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [19:0] tlb_io_tlb_read_port_paddr_1; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [2:0] tlb_io_tlb_read_port_c_0; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire [2:0] tlb_io_tlb_read_port_c_1; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire  tlb_io_tlb_read_port_d_0; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire  tlb_io_tlb_read_port_d_1; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire  tlb_io_tlb_read_port_v_0; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire  tlb_io_tlb_read_port_v_1; // @[double_ports_tlb_for_inst_and_data.scala 49:30]
  wire  tlb_1_clock; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire  tlb_1_reset; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [31:0] tlb_1_io_vaddr; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [31:0] tlb_1_io_paddr; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [7:0] tlb_1_io_cp0_asid; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [3:0] tlb_1_io_tlb_write_index; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [3:0] tlb_1_io_tlb_read_index; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire  tlb_1_io_tlb_write_en; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [3:0] tlb_1_io_tlb_search_index; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire  tlb_1_io_tlb_search_hit; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire  tlb_1_io_tlb_search_ineffective; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire  tlb_1_io_tlb_search_has_changed; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [18:0] tlb_1_io_tlb_write_port_vaddr; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [7:0] tlb_1_io_tlb_write_port_asid; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire  tlb_1_io_tlb_write_port_g; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [19:0] tlb_1_io_tlb_write_port_paddr_0; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [19:0] tlb_1_io_tlb_write_port_paddr_1; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [2:0] tlb_1_io_tlb_write_port_c_0; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [2:0] tlb_1_io_tlb_write_port_c_1; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire  tlb_1_io_tlb_write_port_d_0; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire  tlb_1_io_tlb_write_port_d_1; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire  tlb_1_io_tlb_write_port_v_0; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire  tlb_1_io_tlb_write_port_v_1; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [18:0] tlb_1_io_tlb_read_port_vaddr; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [7:0] tlb_1_io_tlb_read_port_asid; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire  tlb_1_io_tlb_read_port_g; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [19:0] tlb_1_io_tlb_read_port_paddr_0; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [19:0] tlb_1_io_tlb_read_port_paddr_1; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [2:0] tlb_1_io_tlb_read_port_c_0; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire [2:0] tlb_1_io_tlb_read_port_c_1; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire  tlb_1_io_tlb_read_port_d_0; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire  tlb_1_io_tlb_read_port_d_1; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire  tlb_1_io_tlb_read_port_v_0; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  wire  tlb_1_io_tlb_read_port_v_1; // @[double_ports_tlb_for_inst_and_data.scala 50:30]
  tlb tlb ( // @[double_ports_tlb_for_inst_and_data.scala 49:30]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_vaddr(tlb_io_vaddr),
    .io_paddr(tlb_io_paddr),
    .io_cp0_asid(tlb_io_cp0_asid),
    .io_tlb_write_index(tlb_io_tlb_write_index),
    .io_tlb_read_index(tlb_io_tlb_read_index),
    .io_tlb_write_en(tlb_io_tlb_write_en),
    .io_tlb_search_index(tlb_io_tlb_search_index),
    .io_tlb_search_hit(tlb_io_tlb_search_hit),
    .io_tlb_search_ineffective(tlb_io_tlb_search_ineffective),
    .io_tlb_search_has_changed(tlb_io_tlb_search_has_changed),
    .io_tlb_write_port_vaddr(tlb_io_tlb_write_port_vaddr),
    .io_tlb_write_port_asid(tlb_io_tlb_write_port_asid),
    .io_tlb_write_port_g(tlb_io_tlb_write_port_g),
    .io_tlb_write_port_paddr_0(tlb_io_tlb_write_port_paddr_0),
    .io_tlb_write_port_paddr_1(tlb_io_tlb_write_port_paddr_1),
    .io_tlb_write_port_c_0(tlb_io_tlb_write_port_c_0),
    .io_tlb_write_port_c_1(tlb_io_tlb_write_port_c_1),
    .io_tlb_write_port_d_0(tlb_io_tlb_write_port_d_0),
    .io_tlb_write_port_d_1(tlb_io_tlb_write_port_d_1),
    .io_tlb_write_port_v_0(tlb_io_tlb_write_port_v_0),
    .io_tlb_write_port_v_1(tlb_io_tlb_write_port_v_1),
    .io_tlb_read_port_vaddr(tlb_io_tlb_read_port_vaddr),
    .io_tlb_read_port_asid(tlb_io_tlb_read_port_asid),
    .io_tlb_read_port_g(tlb_io_tlb_read_port_g),
    .io_tlb_read_port_paddr_0(tlb_io_tlb_read_port_paddr_0),
    .io_tlb_read_port_paddr_1(tlb_io_tlb_read_port_paddr_1),
    .io_tlb_read_port_c_0(tlb_io_tlb_read_port_c_0),
    .io_tlb_read_port_c_1(tlb_io_tlb_read_port_c_1),
    .io_tlb_read_port_d_0(tlb_io_tlb_read_port_d_0),
    .io_tlb_read_port_d_1(tlb_io_tlb_read_port_d_1),
    .io_tlb_read_port_v_0(tlb_io_tlb_read_port_v_0),
    .io_tlb_read_port_v_1(tlb_io_tlb_read_port_v_1)
  );
  tlb tlb_1 ( // @[double_ports_tlb_for_inst_and_data.scala 50:30]
    .clock(tlb_1_clock),
    .reset(tlb_1_reset),
    .io_vaddr(tlb_1_io_vaddr),
    .io_paddr(tlb_1_io_paddr),
    .io_cp0_asid(tlb_1_io_cp0_asid),
    .io_tlb_write_index(tlb_1_io_tlb_write_index),
    .io_tlb_read_index(tlb_1_io_tlb_read_index),
    .io_tlb_write_en(tlb_1_io_tlb_write_en),
    .io_tlb_search_index(tlb_1_io_tlb_search_index),
    .io_tlb_search_hit(tlb_1_io_tlb_search_hit),
    .io_tlb_search_ineffective(tlb_1_io_tlb_search_ineffective),
    .io_tlb_search_has_changed(tlb_1_io_tlb_search_has_changed),
    .io_tlb_write_port_vaddr(tlb_1_io_tlb_write_port_vaddr),
    .io_tlb_write_port_asid(tlb_1_io_tlb_write_port_asid),
    .io_tlb_write_port_g(tlb_1_io_tlb_write_port_g),
    .io_tlb_write_port_paddr_0(tlb_1_io_tlb_write_port_paddr_0),
    .io_tlb_write_port_paddr_1(tlb_1_io_tlb_write_port_paddr_1),
    .io_tlb_write_port_c_0(tlb_1_io_tlb_write_port_c_0),
    .io_tlb_write_port_c_1(tlb_1_io_tlb_write_port_c_1),
    .io_tlb_write_port_d_0(tlb_1_io_tlb_write_port_d_0),
    .io_tlb_write_port_d_1(tlb_1_io_tlb_write_port_d_1),
    .io_tlb_write_port_v_0(tlb_1_io_tlb_write_port_v_0),
    .io_tlb_write_port_v_1(tlb_1_io_tlb_write_port_v_1),
    .io_tlb_read_port_vaddr(tlb_1_io_tlb_read_port_vaddr),
    .io_tlb_read_port_asid(tlb_1_io_tlb_read_port_asid),
    .io_tlb_read_port_g(tlb_1_io_tlb_read_port_g),
    .io_tlb_read_port_paddr_0(tlb_1_io_tlb_read_port_paddr_0),
    .io_tlb_read_port_paddr_1(tlb_1_io_tlb_read_port_paddr_1),
    .io_tlb_read_port_c_0(tlb_1_io_tlb_read_port_c_0),
    .io_tlb_read_port_c_1(tlb_1_io_tlb_read_port_c_1),
    .io_tlb_read_port_d_0(tlb_1_io_tlb_read_port_d_0),
    .io_tlb_read_port_d_1(tlb_1_io_tlb_read_port_d_1),
    .io_tlb_read_port_v_0(tlb_1_io_tlb_read_port_v_0),
    .io_tlb_read_port_v_1(tlb_1_io_tlb_read_port_v_1)
  );
  assign io_tlb_search_index = tlb_1_io_tlb_search_index; // @[double_ports_tlb_for_inst_and_data.scala 74:25]
  assign io_tlb_search_hit = tlb_1_io_tlb_search_hit; // @[double_ports_tlb_for_inst_and_data.scala 86:23]
  assign io_tlb_dirty_exception = io_dcache_port_wr & tlb_1_io_tlb_search_has_changed & io_dcache_port_req; // @[double_ports_tlb_for_inst_and_data.scala 84:90]
  assign io_tlb_read_port_vaddr = tlb_1_io_tlb_read_port_vaddr; // @[double_ports_tlb_for_inst_and_data.scala 73:22]
  assign io_tlb_read_port_asid = tlb_1_io_tlb_read_port_asid; // @[double_ports_tlb_for_inst_and_data.scala 73:22]
  assign io_tlb_read_port_g = tlb_1_io_tlb_read_port_g; // @[double_ports_tlb_for_inst_and_data.scala 73:22]
  assign io_tlb_read_port_paddr_0 = tlb_1_io_tlb_read_port_paddr_0; // @[double_ports_tlb_for_inst_and_data.scala 73:22]
  assign io_tlb_read_port_paddr_1 = tlb_1_io_tlb_read_port_paddr_1; // @[double_ports_tlb_for_inst_and_data.scala 73:22]
  assign io_tlb_read_port_c_0 = tlb_1_io_tlb_read_port_c_0; // @[double_ports_tlb_for_inst_and_data.scala 73:22]
  assign io_tlb_read_port_c_1 = tlb_1_io_tlb_read_port_c_1; // @[double_ports_tlb_for_inst_and_data.scala 73:22]
  assign io_tlb_read_port_d_0 = tlb_1_io_tlb_read_port_d_0; // @[double_ports_tlb_for_inst_and_data.scala 73:22]
  assign io_tlb_read_port_d_1 = tlb_1_io_tlb_read_port_d_1; // @[double_ports_tlb_for_inst_and_data.scala 73:22]
  assign io_tlb_read_port_v_0 = tlb_1_io_tlb_read_port_v_0; // @[double_ports_tlb_for_inst_and_data.scala 73:22]
  assign io_tlb_read_port_v_1 = tlb_1_io_tlb_read_port_v_1; // @[double_ports_tlb_for_inst_and_data.scala 73:22]
  assign io_icache_port_paddr = tlb_io_paddr; // @[double_ports_tlb_for_inst_and_data.scala 56:26]
  assign io_icache_port_tlb_search_not_hit_exception = ~tlb_io_tlb_search_hit & io_icache_port_req; // @[double_ports_tlb_for_inst_and_data.scala 79:85]
  assign io_icache_port_tlb_search_ineffective_exception = tlb_io_tlb_search_ineffective & io_icache_port_req; // @[double_ports_tlb_for_inst_and_data.scala 78:92]
  assign io_dcache_port_paddr = tlb_1_io_paddr; // @[double_ports_tlb_for_inst_and_data.scala 55:26]
  assign io_dcache_port_tlb_search_not_hit_exception = ~tlb_1_io_tlb_search_hit & io_dcache_port_req; // @[double_ports_tlb_for_inst_and_data.scala 82:85]
  assign io_dcache_port_tlb_search_ineffective_exception = tlb_1_io_tlb_search_ineffective & io_dcache_port_req; // @[double_ports_tlb_for_inst_and_data.scala 81:92]
  assign tlb_clock = clock;
  assign tlb_reset = reset;
  assign tlb_io_vaddr = io_icache_port_vaddr; // @[double_ports_tlb_for_inst_and_data.scala 52:24]
  assign tlb_io_cp0_asid = io_cp0_asid; // @[double_ports_tlb_for_inst_and_data.scala 64:34]
  assign tlb_io_tlb_write_index = io_tlb_write_index; // @[double_ports_tlb_for_inst_and_data.scala 63:34]
  assign tlb_io_tlb_read_index = 4'h0; // @[double_ports_tlb_for_inst_and_data.scala 65:34]
  assign tlb_io_tlb_write_en = io_tlb_write_en; // @[double_ports_tlb_for_inst_and_data.scala 62:34]
  assign tlb_io_tlb_write_port_vaddr = io_tlb_write_port_vaddr; // @[double_ports_tlb_for_inst_and_data.scala 61:34]
  assign tlb_io_tlb_write_port_asid = io_tlb_write_port_asid; // @[double_ports_tlb_for_inst_and_data.scala 61:34]
  assign tlb_io_tlb_write_port_g = io_tlb_write_port_g; // @[double_ports_tlb_for_inst_and_data.scala 61:34]
  assign tlb_io_tlb_write_port_paddr_0 = io_tlb_write_port_paddr_0; // @[double_ports_tlb_for_inst_and_data.scala 61:34]
  assign tlb_io_tlb_write_port_paddr_1 = io_tlb_write_port_paddr_1; // @[double_ports_tlb_for_inst_and_data.scala 61:34]
  assign tlb_io_tlb_write_port_c_0 = io_tlb_write_port_c_0; // @[double_ports_tlb_for_inst_and_data.scala 61:34]
  assign tlb_io_tlb_write_port_c_1 = io_tlb_write_port_c_1; // @[double_ports_tlb_for_inst_and_data.scala 61:34]
  assign tlb_io_tlb_write_port_d_0 = io_tlb_write_port_d_0; // @[double_ports_tlb_for_inst_and_data.scala 61:34]
  assign tlb_io_tlb_write_port_d_1 = io_tlb_write_port_d_1; // @[double_ports_tlb_for_inst_and_data.scala 61:34]
  assign tlb_io_tlb_write_port_v_0 = io_tlb_write_port_v_0; // @[double_ports_tlb_for_inst_and_data.scala 61:34]
  assign tlb_io_tlb_write_port_v_1 = io_tlb_write_port_v_1; // @[double_ports_tlb_for_inst_and_data.scala 61:34]
  assign tlb_1_clock = clock;
  assign tlb_1_reset = reset;
  assign tlb_1_io_vaddr = io_dcache_port_vaddr; // @[double_ports_tlb_for_inst_and_data.scala 53:24]
  assign tlb_1_io_cp0_asid = io_cp0_asid; // @[double_ports_tlb_for_inst_and_data.scala 71:34]
  assign tlb_1_io_tlb_write_index = io_tlb_write_index; // @[double_ports_tlb_for_inst_and_data.scala 70:34]
  assign tlb_1_io_tlb_read_index = io_tlb_read_index; // @[double_ports_tlb_for_inst_and_data.scala 72:34]
  assign tlb_1_io_tlb_write_en = io_tlb_write_en; // @[double_ports_tlb_for_inst_and_data.scala 69:34]
  assign tlb_1_io_tlb_write_port_vaddr = io_tlb_write_port_vaddr; // @[double_ports_tlb_for_inst_and_data.scala 68:34]
  assign tlb_1_io_tlb_write_port_asid = io_tlb_write_port_asid; // @[double_ports_tlb_for_inst_and_data.scala 68:34]
  assign tlb_1_io_tlb_write_port_g = io_tlb_write_port_g; // @[double_ports_tlb_for_inst_and_data.scala 68:34]
  assign tlb_1_io_tlb_write_port_paddr_0 = io_tlb_write_port_paddr_0; // @[double_ports_tlb_for_inst_and_data.scala 68:34]
  assign tlb_1_io_tlb_write_port_paddr_1 = io_tlb_write_port_paddr_1; // @[double_ports_tlb_for_inst_and_data.scala 68:34]
  assign tlb_1_io_tlb_write_port_c_0 = io_tlb_write_port_c_0; // @[double_ports_tlb_for_inst_and_data.scala 68:34]
  assign tlb_1_io_tlb_write_port_c_1 = io_tlb_write_port_c_1; // @[double_ports_tlb_for_inst_and_data.scala 68:34]
  assign tlb_1_io_tlb_write_port_d_0 = io_tlb_write_port_d_0; // @[double_ports_tlb_for_inst_and_data.scala 68:34]
  assign tlb_1_io_tlb_write_port_d_1 = io_tlb_write_port_d_1; // @[double_ports_tlb_for_inst_and_data.scala 68:34]
  assign tlb_1_io_tlb_write_port_v_0 = io_tlb_write_port_v_0; // @[double_ports_tlb_for_inst_and_data.scala 68:34]
  assign tlb_1_io_tlb_write_port_v_1 = io_tlb_write_port_v_1; // @[double_ports_tlb_for_inst_and_data.scala 68:34]
endmodule
module mycpu_top(
  input         aresetn,
  input         aclk,
  input  [5:0]  ext_int,
  output [3:0]  arid,
  output [31:0] araddr,
  output [3:0]  arlen,
  output [2:0]  arsize,
  output [1:0]  arburst,
  output [1:0]  arlock,
  output [3:0]  arcache,
  output [2:0]  arprot,
  output        arvalid,
  input         arready,
  input  [3:0]  rid,
  input  [31:0] rdata,
  input  [1:0]  rresp,
  input         rlast,
  input         rvalid,
  output        rready,
  output [3:0]  awid,
  output [31:0] awaddr,
  output [3:0]  awlen,
  output [2:0]  awsize,
  output [1:0]  awburst,
  output [1:0]  awlock,
  output [3:0]  awcache,
  output [2:0]  awprot,
  output        awvalid,
  input         awready,
  output [3:0]  wid,
  output [31:0] wdata,
  output [3:0]  wstrb,
  output        wlast,
  output        wvalid,
  input         wready,
  input  [3:0]  bid,
  input  [1:0]  bresp,
  input         bvalid,
  output        bready,
  output [31:0] debug_wb_pc,
  output [3:0]  debug_wb_rf_wen,
  output [4:0]  debug_wb_rf_wnum,
  output [31:0] debug_wb_rf_wdata
);
  wire  u_axi_cache_bridge_aclk; // @[my_cpu_top.scala 318:36]
  wire  u_axi_cache_bridge_aresetn; // @[my_cpu_top.scala 318:36]
  wire [7:0] u_axi_cache_bridge_s_axi_awid; // @[my_cpu_top.scala 318:36]
  wire [63:0] u_axi_cache_bridge_s_axi_awaddr; // @[my_cpu_top.scala 318:36]
  wire [7:0] u_axi_cache_bridge_s_axi_awlen; // @[my_cpu_top.scala 318:36]
  wire [5:0] u_axi_cache_bridge_s_axi_awsize; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_s_axi_awburst; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_s_axi_awlock; // @[my_cpu_top.scala 318:36]
  wire [7:0] u_axi_cache_bridge_s_axi_awcache; // @[my_cpu_top.scala 318:36]
  wire [5:0] u_axi_cache_bridge_s_axi_awprot; // @[my_cpu_top.scala 318:36]
  wire [7:0] u_axi_cache_bridge_s_axi_awqos; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_s_axi_awvalid; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_s_axi_awready; // @[my_cpu_top.scala 318:36]
  wire [7:0] u_axi_cache_bridge_s_axi_wid; // @[my_cpu_top.scala 318:36]
  wire [63:0] u_axi_cache_bridge_s_axi_wdata; // @[my_cpu_top.scala 318:36]
  wire [7:0] u_axi_cache_bridge_s_axi_wstrb; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_s_axi_wlast; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_s_axi_wvalid; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_s_axi_wready; // @[my_cpu_top.scala 318:36]
  wire [7:0] u_axi_cache_bridge_s_axi_bid; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_s_axi_bresp; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_s_axi_bvalid; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_s_axi_bready; // @[my_cpu_top.scala 318:36]
  wire [7:0] u_axi_cache_bridge_s_axi_arid; // @[my_cpu_top.scala 318:36]
  wire [63:0] u_axi_cache_bridge_s_axi_araddr; // @[my_cpu_top.scala 318:36]
  wire [7:0] u_axi_cache_bridge_s_axi_arlen; // @[my_cpu_top.scala 318:36]
  wire [5:0] u_axi_cache_bridge_s_axi_arsize; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_s_axi_arburst; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_s_axi_arlock; // @[my_cpu_top.scala 318:36]
  wire [7:0] u_axi_cache_bridge_s_axi_arcache; // @[my_cpu_top.scala 318:36]
  wire [5:0] u_axi_cache_bridge_s_axi_arprot; // @[my_cpu_top.scala 318:36]
  wire [7:0] u_axi_cache_bridge_s_axi_arqos; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_s_axi_arvalid; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_s_axi_arready; // @[my_cpu_top.scala 318:36]
  wire [7:0] u_axi_cache_bridge_s_axi_rid; // @[my_cpu_top.scala 318:36]
  wire [63:0] u_axi_cache_bridge_s_axi_rdata; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_s_axi_rresp; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_s_axi_rlast; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_s_axi_rvalid; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_s_axi_rready; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_m_axi_awid; // @[my_cpu_top.scala 318:36]
  wire [31:0] u_axi_cache_bridge_m_axi_awaddr; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_m_axi_awlen; // @[my_cpu_top.scala 318:36]
  wire [2:0] u_axi_cache_bridge_m_axi_awsize; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_m_axi_awburst; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_m_axi_awlock; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_m_axi_awcache; // @[my_cpu_top.scala 318:36]
  wire [2:0] u_axi_cache_bridge_m_axi_awprot; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_m_axi_awqos; // @[my_cpu_top.scala 318:36]
  wire  u_axi_cache_bridge_m_axi_awvalid; // @[my_cpu_top.scala 318:36]
  wire  u_axi_cache_bridge_m_axi_awready; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_m_axi_wid; // @[my_cpu_top.scala 318:36]
  wire [31:0] u_axi_cache_bridge_m_axi_wdata; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_m_axi_wstrb; // @[my_cpu_top.scala 318:36]
  wire  u_axi_cache_bridge_m_axi_wlast; // @[my_cpu_top.scala 318:36]
  wire  u_axi_cache_bridge_m_axi_wvalid; // @[my_cpu_top.scala 318:36]
  wire  u_axi_cache_bridge_m_axi_wready; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_m_axi_bid; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_m_axi_bresp; // @[my_cpu_top.scala 318:36]
  wire  u_axi_cache_bridge_m_axi_bvalid; // @[my_cpu_top.scala 318:36]
  wire  u_axi_cache_bridge_m_axi_bready; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_m_axi_arid; // @[my_cpu_top.scala 318:36]
  wire [31:0] u_axi_cache_bridge_m_axi_araddr; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_m_axi_arlen; // @[my_cpu_top.scala 318:36]
  wire [2:0] u_axi_cache_bridge_m_axi_arsize; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_m_axi_arburst; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_m_axi_arlock; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_m_axi_arcache; // @[my_cpu_top.scala 318:36]
  wire [2:0] u_axi_cache_bridge_m_axi_arprot; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_m_axi_arqos; // @[my_cpu_top.scala 318:36]
  wire  u_axi_cache_bridge_m_axi_arvalid; // @[my_cpu_top.scala 318:36]
  wire  u_axi_cache_bridge_m_axi_rready; // @[my_cpu_top.scala 318:36]
  wire  u_axi_cache_bridge_m_axi_arready; // @[my_cpu_top.scala 318:36]
  wire [3:0] u_axi_cache_bridge_m_axi_rid; // @[my_cpu_top.scala 318:36]
  wire [31:0] u_axi_cache_bridge_m_axi_rdata; // @[my_cpu_top.scala 318:36]
  wire [1:0] u_axi_cache_bridge_m_axi_rresp; // @[my_cpu_top.scala 318:36]
  wire  u_axi_cache_bridge_m_axi_rlast; // @[my_cpu_top.scala 318:36]
  wire  u_axi_cache_bridge_m_axi_rvalid; // @[my_cpu_top.scala 318:36]
  wire [5:0] u_mips_cpu_ext_int; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_resetn; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_clk; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_inst_cache; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_inst_sram_en; // @[my_cpu_top.scala 319:28]
  wire [31:0] u_mips_cpu_inst_sram_addr; // @[my_cpu_top.scala 319:28]
  wire [39:0] u_mips_cpu_inst_sram_rdata_L; // @[my_cpu_top.scala 319:28]
  wire [1:0] u_mips_cpu_inst_write_en; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_inst_ready_branch; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_inst_buffer_empty; // @[my_cpu_top.scala 319:28]
  wire [7:0] u_mips_cpu_cp0_asid; // @[my_cpu_top.scala 319:28]
  wire [1:0] u_mips_cpu_inst_tlb_exception; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_stage2_flush; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_stage2_stall; // @[my_cpu_top.scala 319:28]
  wire [1:0] u_mips_cpu_stage1_valid_flush; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_inst_ready_to_use; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_inst_buffer_full; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_data_sram_en; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_data_sram_wen; // @[my_cpu_top.scala 319:28]
  wire [1:0] u_mips_cpu_data_size; // @[my_cpu_top.scala 319:28]
  wire [31:0] u_mips_cpu_data_sram_addr; // @[my_cpu_top.scala 319:28]
  wire [31:0] u_mips_cpu_data_sram_wdata; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_data_cache; // @[my_cpu_top.scala 319:28]
  wire [31:0] u_mips_cpu_data_sram_rdata; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_data_stage2_stall; // @[my_cpu_top.scala 319:28]
  wire [2:0] u_mips_cpu_data_tlb_exception; // @[my_cpu_top.scala 319:28]
  wire [3:0] u_mips_cpu_data_wstrb; // @[my_cpu_top.scala 319:28]
  wire [31:0] u_mips_cpu_tlbp_search_vaddr; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_tlbp_search_en; // @[my_cpu_top.scala 319:28]
  wire [3:0] u_mips_cpu_tlb_search_index; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_tlb_search_hit; // @[my_cpu_top.scala 319:28]
  wire [3:0] u_mips_cpu_tlb_read_index; // @[my_cpu_top.scala 319:28]
  wire [3:0] u_mips_cpu_tlb_write_index; // @[my_cpu_top.scala 319:28]
  wire [31:0] u_mips_cpu_debug_wb_pc; // @[my_cpu_top.scala 319:28]
  wire [3:0] u_mips_cpu_debug_wb_rf_wen; // @[my_cpu_top.scala 319:28]
  wire [4:0] u_mips_cpu_debug_wb_rf_wnum; // @[my_cpu_top.scala 319:28]
  wire [31:0] u_mips_cpu_debug_wb_rf_wdata; // @[my_cpu_top.scala 319:28]
  wire [18:0] u_mips_cpu_cp0_tlb_read_data_vaddr; // @[my_cpu_top.scala 319:28]
  wire [7:0] u_mips_cpu_cp0_tlb_read_data_asid; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_cp0_tlb_read_data_g; // @[my_cpu_top.scala 319:28]
  wire [19:0] u_mips_cpu_cp0_tlb_read_data_paddr_0; // @[my_cpu_top.scala 319:28]
  wire [19:0] u_mips_cpu_cp0_tlb_read_data_paddr_1; // @[my_cpu_top.scala 319:28]
  wire [2:0] u_mips_cpu_cp0_tlb_read_data_c_0; // @[my_cpu_top.scala 319:28]
  wire [2:0] u_mips_cpu_cp0_tlb_read_data_c_1; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_cp0_tlb_read_data_d_0; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_cp0_tlb_read_data_d_1; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_cp0_tlb_read_data_v_0; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_cp0_tlb_read_data_v_1; // @[my_cpu_top.scala 319:28]
  wire [18:0] u_mips_cpu_cp0_tlb_write_data_vaddr; // @[my_cpu_top.scala 319:28]
  wire [7:0] u_mips_cpu_cp0_tlb_write_data_asid; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_cp0_tlb_write_data_g; // @[my_cpu_top.scala 319:28]
  wire [19:0] u_mips_cpu_cp0_tlb_write_data_paddr_0; // @[my_cpu_top.scala 319:28]
  wire [19:0] u_mips_cpu_cp0_tlb_write_data_paddr_1; // @[my_cpu_top.scala 319:28]
  wire [2:0] u_mips_cpu_cp0_tlb_write_data_c_0; // @[my_cpu_top.scala 319:28]
  wire [2:0] u_mips_cpu_cp0_tlb_write_data_c_1; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_cp0_tlb_write_data_d_0; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_cp0_tlb_write_data_d_1; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_cp0_tlb_write_data_v_0; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_cp0_tlb_write_data_v_1; // @[my_cpu_top.scala 319:28]
  wire  u_mips_cpu_tlb_write_en; // @[my_cpu_top.scala 319:28]
  wire  inst_cache_clock; // @[my_cpu_top.scala 320:30]
  wire  inst_cache_reset; // @[my_cpu_top.scala 320:30]
  wire [31:0] inst_cache_io_port_araddr; // @[my_cpu_top.scala 320:30]
  wire [3:0] inst_cache_io_port_arlen; // @[my_cpu_top.scala 320:30]
  wire [1:0] inst_cache_io_port_arburst; // @[my_cpu_top.scala 320:30]
  wire  inst_cache_io_port_arvalid; // @[my_cpu_top.scala 320:30]
  wire  inst_cache_io_port_arready; // @[my_cpu_top.scala 320:30]
  wire [31:0] inst_cache_io_port_rdata; // @[my_cpu_top.scala 320:30]
  wire  inst_cache_io_port_rlast; // @[my_cpu_top.scala 320:30]
  wire  inst_cache_io_port_rvalid; // @[my_cpu_top.scala 320:30]
  wire  inst_cache_io_port_sram_req; // @[my_cpu_top.scala 320:30]
  wire [31:0] inst_cache_io_port_sram_addr; // @[my_cpu_top.scala 320:30]
  wire [1:0] inst_cache_io_port_sram_write_en; // @[my_cpu_top.scala 320:30]
  wire [39:0] inst_cache_io_port_sram_rdata_L; // @[my_cpu_top.scala 320:30]
  wire  inst_cache_io_port_sram_cache; // @[my_cpu_top.scala 320:30]
  wire  inst_cache_io_stage2_flush; // @[my_cpu_top.scala 320:30]
  wire  inst_cache_io_stage2_stall; // @[my_cpu_top.scala 320:30]
  wire [1:0] inst_cache_io_stage1_valid_flush; // @[my_cpu_top.scala 320:30]
  wire  inst_cache_io_inst_ready_to_use; // @[my_cpu_top.scala 320:30]
  wire  inst_cache_io_inst_buffer_full; // @[my_cpu_top.scala 320:30]
  wire [1:0] inst_cache_io_stage2_exception; // @[my_cpu_top.scala 320:30]
  wire [7:0] inst_cache_io_cp0_asid; // @[my_cpu_top.scala 320:30]
  wire [31:0] inst_cache_io_v_addr_for_tlb; // @[my_cpu_top.scala 320:30]
  wire [31:0] inst_cache_io_p_addr_for_tlb; // @[my_cpu_top.scala 320:30]
  wire  inst_cache_io_tlb_req; // @[my_cpu_top.scala 320:30]
  wire [1:0] inst_cache_io_tlb_exception; // @[my_cpu_top.scala 320:30]
  wire  inst_cache_io_inst_ready_branch; // @[my_cpu_top.scala 320:30]
  wire  inst_cache_io_inst_buffer_empty; // @[my_cpu_top.scala 320:30]
  wire  data_cache_clock; // @[my_cpu_top.scala 322:30]
  wire  data_cache_reset; // @[my_cpu_top.scala 322:30]
  wire [31:0] data_cache_io_port_araddr; // @[my_cpu_top.scala 322:30]
  wire [3:0] data_cache_io_port_arlen; // @[my_cpu_top.scala 322:30]
  wire [2:0] data_cache_io_port_arsize; // @[my_cpu_top.scala 322:30]
  wire [1:0] data_cache_io_port_arburst; // @[my_cpu_top.scala 322:30]
  wire  data_cache_io_port_arvalid; // @[my_cpu_top.scala 322:30]
  wire  data_cache_io_port_arready; // @[my_cpu_top.scala 322:30]
  wire [31:0] data_cache_io_port_rdata; // @[my_cpu_top.scala 322:30]
  wire  data_cache_io_port_rlast; // @[my_cpu_top.scala 322:30]
  wire  data_cache_io_port_rvalid; // @[my_cpu_top.scala 322:30]
  wire [31:0] data_cache_io_port_awaddr; // @[my_cpu_top.scala 322:30]
  wire [3:0] data_cache_io_port_awlen; // @[my_cpu_top.scala 322:30]
  wire [2:0] data_cache_io_port_awsize; // @[my_cpu_top.scala 322:30]
  wire [1:0] data_cache_io_port_awburst; // @[my_cpu_top.scala 322:30]
  wire  data_cache_io_port_awvalid; // @[my_cpu_top.scala 322:30]
  wire  data_cache_io_port_awready; // @[my_cpu_top.scala 322:30]
  wire [31:0] data_cache_io_port_wdata; // @[my_cpu_top.scala 322:30]
  wire [3:0] data_cache_io_port_wstrb; // @[my_cpu_top.scala 322:30]
  wire  data_cache_io_port_wlast; // @[my_cpu_top.scala 322:30]
  wire  data_cache_io_port_wvalid; // @[my_cpu_top.scala 322:30]
  wire  data_cache_io_port_wready; // @[my_cpu_top.scala 322:30]
  wire  data_cache_io_port_bvalid; // @[my_cpu_top.scala 322:30]
  wire  data_cache_io_port_sram_req; // @[my_cpu_top.scala 322:30]
  wire  data_cache_io_port_sram_wr; // @[my_cpu_top.scala 322:30]
  wire [1:0] data_cache_io_port_sram_size; // @[my_cpu_top.scala 322:30]
  wire [31:0] data_cache_io_port_sram_addr; // @[my_cpu_top.scala 322:30]
  wire [31:0] data_cache_io_port_sram_wdata; // @[my_cpu_top.scala 322:30]
  wire [31:0] data_cache_io_port_sram_rdata; // @[my_cpu_top.scala 322:30]
  wire  data_cache_io_port_sram_cache; // @[my_cpu_top.scala 322:30]
  wire  data_cache_io_stage2_stall; // @[my_cpu_top.scala 322:30]
  wire  data_cache_io_stage1_wr; // @[my_cpu_top.scala 322:30]
  wire [31:0] data_cache_io_v_addr_for_tlb; // @[my_cpu_top.scala 322:30]
  wire [31:0] data_cache_io_p_addr_for_tlb; // @[my_cpu_top.scala 322:30]
  wire  data_cache_io_tlb_req; // @[my_cpu_top.scala 322:30]
  wire [2:0] data_cache_io_tlb_exception; // @[my_cpu_top.scala 322:30]
  wire [2:0] data_cache_io_stage1_tlb_exception; // @[my_cpu_top.scala 322:30]
  wire [3:0] data_cache_io_data_wstrb; // @[my_cpu_top.scala 322:30]
  wire  double_ports_tlb_for_inst_and_data_clock; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_reset; // @[my_cpu_top.scala 325:22]
  wire [7:0] double_ports_tlb_for_inst_and_data_io_cp0_asid; // @[my_cpu_top.scala 325:22]
  wire [3:0] double_ports_tlb_for_inst_and_data_io_tlb_write_index; // @[my_cpu_top.scala 325:22]
  wire [3:0] double_ports_tlb_for_inst_and_data_io_tlb_read_index; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_tlb_write_en; // @[my_cpu_top.scala 325:22]
  wire [3:0] double_ports_tlb_for_inst_and_data_io_tlb_search_index; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_tlb_search_hit; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_tlb_dirty_exception; // @[my_cpu_top.scala 325:22]
  wire [18:0] double_ports_tlb_for_inst_and_data_io_tlb_write_port_vaddr; // @[my_cpu_top.scala 325:22]
  wire [7:0] double_ports_tlb_for_inst_and_data_io_tlb_write_port_asid; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_tlb_write_port_g; // @[my_cpu_top.scala 325:22]
  wire [19:0] double_ports_tlb_for_inst_and_data_io_tlb_write_port_paddr_0; // @[my_cpu_top.scala 325:22]
  wire [19:0] double_ports_tlb_for_inst_and_data_io_tlb_write_port_paddr_1; // @[my_cpu_top.scala 325:22]
  wire [2:0] double_ports_tlb_for_inst_and_data_io_tlb_write_port_c_0; // @[my_cpu_top.scala 325:22]
  wire [2:0] double_ports_tlb_for_inst_and_data_io_tlb_write_port_c_1; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_tlb_write_port_d_0; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_tlb_write_port_d_1; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_tlb_write_port_v_0; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_tlb_write_port_v_1; // @[my_cpu_top.scala 325:22]
  wire [18:0] double_ports_tlb_for_inst_and_data_io_tlb_read_port_vaddr; // @[my_cpu_top.scala 325:22]
  wire [7:0] double_ports_tlb_for_inst_and_data_io_tlb_read_port_asid; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_tlb_read_port_g; // @[my_cpu_top.scala 325:22]
  wire [19:0] double_ports_tlb_for_inst_and_data_io_tlb_read_port_paddr_0; // @[my_cpu_top.scala 325:22]
  wire [19:0] double_ports_tlb_for_inst_and_data_io_tlb_read_port_paddr_1; // @[my_cpu_top.scala 325:22]
  wire [2:0] double_ports_tlb_for_inst_and_data_io_tlb_read_port_c_0; // @[my_cpu_top.scala 325:22]
  wire [2:0] double_ports_tlb_for_inst_and_data_io_tlb_read_port_c_1; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_tlb_read_port_d_0; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_tlb_read_port_d_1; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_tlb_read_port_v_0; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_tlb_read_port_v_1; // @[my_cpu_top.scala 325:22]
  wire [31:0] double_ports_tlb_for_inst_and_data_io_icache_port_vaddr; // @[my_cpu_top.scala 325:22]
  wire [31:0] double_ports_tlb_for_inst_and_data_io_icache_port_paddr; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_icache_port_req; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_icache_port_tlb_search_not_hit_exception; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_icache_port_tlb_search_ineffective_exception; // @[my_cpu_top.scala 325:22]
  wire [31:0] double_ports_tlb_for_inst_and_data_io_dcache_port_vaddr; // @[my_cpu_top.scala 325:22]
  wire [31:0] double_ports_tlb_for_inst_and_data_io_dcache_port_paddr; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_dcache_port_req; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_dcache_port_wr; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_dcache_port_tlb_search_not_hit_exception; // @[my_cpu_top.scala 325:22]
  wire  double_ports_tlb_for_inst_and_data_io_dcache_port_tlb_search_ineffective_exception; // @[my_cpu_top.scala 325:22]
  wire [1:0] hi = {double_ports_tlb_for_inst_and_data_io_tlb_dirty_exception,
    double_ports_tlb_for_inst_and_data_io_dcache_port_tlb_search_ineffective_exception}; // @[Cat.scala 31:58]
  axi_crossbar_0 u_axi_cache_bridge ( // @[my_cpu_top.scala 318:36]
    .aclk(u_axi_cache_bridge_aclk),
    .aresetn(u_axi_cache_bridge_aresetn),
    .s_axi_awid(u_axi_cache_bridge_s_axi_awid),
    .s_axi_awaddr(u_axi_cache_bridge_s_axi_awaddr),
    .s_axi_awlen(u_axi_cache_bridge_s_axi_awlen),
    .s_axi_awsize(u_axi_cache_bridge_s_axi_awsize),
    .s_axi_awburst(u_axi_cache_bridge_s_axi_awburst),
    .s_axi_awlock(u_axi_cache_bridge_s_axi_awlock),
    .s_axi_awcache(u_axi_cache_bridge_s_axi_awcache),
    .s_axi_awprot(u_axi_cache_bridge_s_axi_awprot),
    .s_axi_awqos(u_axi_cache_bridge_s_axi_awqos),
    .s_axi_awvalid(u_axi_cache_bridge_s_axi_awvalid),
    .s_axi_awready(u_axi_cache_bridge_s_axi_awready),
    .s_axi_wid(u_axi_cache_bridge_s_axi_wid),
    .s_axi_wdata(u_axi_cache_bridge_s_axi_wdata),
    .s_axi_wstrb(u_axi_cache_bridge_s_axi_wstrb),
    .s_axi_wlast(u_axi_cache_bridge_s_axi_wlast),
    .s_axi_wvalid(u_axi_cache_bridge_s_axi_wvalid),
    .s_axi_wready(u_axi_cache_bridge_s_axi_wready),
    .s_axi_bid(u_axi_cache_bridge_s_axi_bid),
    .s_axi_bresp(u_axi_cache_bridge_s_axi_bresp),
    .s_axi_bvalid(u_axi_cache_bridge_s_axi_bvalid),
    .s_axi_bready(u_axi_cache_bridge_s_axi_bready),
    .s_axi_arid(u_axi_cache_bridge_s_axi_arid),
    .s_axi_araddr(u_axi_cache_bridge_s_axi_araddr),
    .s_axi_arlen(u_axi_cache_bridge_s_axi_arlen),
    .s_axi_arsize(u_axi_cache_bridge_s_axi_arsize),
    .s_axi_arburst(u_axi_cache_bridge_s_axi_arburst),
    .s_axi_arlock(u_axi_cache_bridge_s_axi_arlock),
    .s_axi_arcache(u_axi_cache_bridge_s_axi_arcache),
    .s_axi_arprot(u_axi_cache_bridge_s_axi_arprot),
    .s_axi_arqos(u_axi_cache_bridge_s_axi_arqos),
    .s_axi_arvalid(u_axi_cache_bridge_s_axi_arvalid),
    .s_axi_arready(u_axi_cache_bridge_s_axi_arready),
    .s_axi_rid(u_axi_cache_bridge_s_axi_rid),
    .s_axi_rdata(u_axi_cache_bridge_s_axi_rdata),
    .s_axi_rresp(u_axi_cache_bridge_s_axi_rresp),
    .s_axi_rlast(u_axi_cache_bridge_s_axi_rlast),
    .s_axi_rvalid(u_axi_cache_bridge_s_axi_rvalid),
    .s_axi_rready(u_axi_cache_bridge_s_axi_rready),
    .m_axi_awid(u_axi_cache_bridge_m_axi_awid),
    .m_axi_awaddr(u_axi_cache_bridge_m_axi_awaddr),
    .m_axi_awlen(u_axi_cache_bridge_m_axi_awlen),
    .m_axi_awsize(u_axi_cache_bridge_m_axi_awsize),
    .m_axi_awburst(u_axi_cache_bridge_m_axi_awburst),
    .m_axi_awlock(u_axi_cache_bridge_m_axi_awlock),
    .m_axi_awcache(u_axi_cache_bridge_m_axi_awcache),
    .m_axi_awprot(u_axi_cache_bridge_m_axi_awprot),
    .m_axi_awqos(u_axi_cache_bridge_m_axi_awqos),
    .m_axi_awvalid(u_axi_cache_bridge_m_axi_awvalid),
    .m_axi_awready(u_axi_cache_bridge_m_axi_awready),
    .m_axi_wid(u_axi_cache_bridge_m_axi_wid),
    .m_axi_wdata(u_axi_cache_bridge_m_axi_wdata),
    .m_axi_wstrb(u_axi_cache_bridge_m_axi_wstrb),
    .m_axi_wlast(u_axi_cache_bridge_m_axi_wlast),
    .m_axi_wvalid(u_axi_cache_bridge_m_axi_wvalid),
    .m_axi_wready(u_axi_cache_bridge_m_axi_wready),
    .m_axi_bid(u_axi_cache_bridge_m_axi_bid),
    .m_axi_bresp(u_axi_cache_bridge_m_axi_bresp),
    .m_axi_bvalid(u_axi_cache_bridge_m_axi_bvalid),
    .m_axi_bready(u_axi_cache_bridge_m_axi_bready),
    .m_axi_arid(u_axi_cache_bridge_m_axi_arid),
    .m_axi_araddr(u_axi_cache_bridge_m_axi_araddr),
    .m_axi_arlen(u_axi_cache_bridge_m_axi_arlen),
    .m_axi_arsize(u_axi_cache_bridge_m_axi_arsize),
    .m_axi_arburst(u_axi_cache_bridge_m_axi_arburst),
    .m_axi_arlock(u_axi_cache_bridge_m_axi_arlock),
    .m_axi_arcache(u_axi_cache_bridge_m_axi_arcache),
    .m_axi_arprot(u_axi_cache_bridge_m_axi_arprot),
    .m_axi_arqos(u_axi_cache_bridge_m_axi_arqos),
    .m_axi_arvalid(u_axi_cache_bridge_m_axi_arvalid),
    .m_axi_rready(u_axi_cache_bridge_m_axi_rready),
    .m_axi_arready(u_axi_cache_bridge_m_axi_arready),
    .m_axi_rid(u_axi_cache_bridge_m_axi_rid),
    .m_axi_rdata(u_axi_cache_bridge_m_axi_rdata),
    .m_axi_rresp(u_axi_cache_bridge_m_axi_rresp),
    .m_axi_rlast(u_axi_cache_bridge_m_axi_rlast),
    .m_axi_rvalid(u_axi_cache_bridge_m_axi_rvalid)
  );
  myCPU u_mips_cpu ( // @[my_cpu_top.scala 319:28]
    .ext_int(u_mips_cpu_ext_int),
    .resetn(u_mips_cpu_resetn),
    .clk(u_mips_cpu_clk),
    .inst_cache(u_mips_cpu_inst_cache),
    .inst_sram_en(u_mips_cpu_inst_sram_en),
    .inst_sram_addr(u_mips_cpu_inst_sram_addr),
    .inst_sram_rdata_L(u_mips_cpu_inst_sram_rdata_L),
    .inst_write_en(u_mips_cpu_inst_write_en),
    .inst_ready_branch(u_mips_cpu_inst_ready_branch),
    .inst_buffer_empty(u_mips_cpu_inst_buffer_empty),
    .cp0_asid(u_mips_cpu_cp0_asid),
    .inst_tlb_exception(u_mips_cpu_inst_tlb_exception),
    .stage2_flush(u_mips_cpu_stage2_flush),
    .stage2_stall(u_mips_cpu_stage2_stall),
    .stage1_valid_flush(u_mips_cpu_stage1_valid_flush),
    .inst_ready_to_use(u_mips_cpu_inst_ready_to_use),
    .inst_buffer_full(u_mips_cpu_inst_buffer_full),
    .data_sram_en(u_mips_cpu_data_sram_en),
    .data_sram_wen(u_mips_cpu_data_sram_wen),
    .data_size(u_mips_cpu_data_size),
    .data_sram_addr(u_mips_cpu_data_sram_addr),
    .data_sram_wdata(u_mips_cpu_data_sram_wdata),
    .data_cache(u_mips_cpu_data_cache),
    .data_sram_rdata(u_mips_cpu_data_sram_rdata),
    .data_stage2_stall(u_mips_cpu_data_stage2_stall),
    .data_tlb_exception(u_mips_cpu_data_tlb_exception),
    .data_wstrb(u_mips_cpu_data_wstrb),
    .tlbp_search_vaddr(u_mips_cpu_tlbp_search_vaddr),
    .tlbp_search_en(u_mips_cpu_tlbp_search_en),
    .tlb_search_index(u_mips_cpu_tlb_search_index),
    .tlb_search_hit(u_mips_cpu_tlb_search_hit),
    .tlb_read_index(u_mips_cpu_tlb_read_index),
    .tlb_write_index(u_mips_cpu_tlb_write_index),
    .debug_wb_pc(u_mips_cpu_debug_wb_pc),
    .debug_wb_rf_wen(u_mips_cpu_debug_wb_rf_wen),
    .debug_wb_rf_wnum(u_mips_cpu_debug_wb_rf_wnum),
    .debug_wb_rf_wdata(u_mips_cpu_debug_wb_rf_wdata),
    .cp0_tlb_read_data_vaddr(u_mips_cpu_cp0_tlb_read_data_vaddr),
    .cp0_tlb_read_data_asid(u_mips_cpu_cp0_tlb_read_data_asid),
    .cp0_tlb_read_data_g(u_mips_cpu_cp0_tlb_read_data_g),
    .cp0_tlb_read_data_paddr_0(u_mips_cpu_cp0_tlb_read_data_paddr_0),
    .cp0_tlb_read_data_paddr_1(u_mips_cpu_cp0_tlb_read_data_paddr_1),
    .cp0_tlb_read_data_c_0(u_mips_cpu_cp0_tlb_read_data_c_0),
    .cp0_tlb_read_data_c_1(u_mips_cpu_cp0_tlb_read_data_c_1),
    .cp0_tlb_read_data_d_0(u_mips_cpu_cp0_tlb_read_data_d_0),
    .cp0_tlb_read_data_d_1(u_mips_cpu_cp0_tlb_read_data_d_1),
    .cp0_tlb_read_data_v_0(u_mips_cpu_cp0_tlb_read_data_v_0),
    .cp0_tlb_read_data_v_1(u_mips_cpu_cp0_tlb_read_data_v_1),
    .cp0_tlb_write_data_vaddr(u_mips_cpu_cp0_tlb_write_data_vaddr),
    .cp0_tlb_write_data_asid(u_mips_cpu_cp0_tlb_write_data_asid),
    .cp0_tlb_write_data_g(u_mips_cpu_cp0_tlb_write_data_g),
    .cp0_tlb_write_data_paddr_0(u_mips_cpu_cp0_tlb_write_data_paddr_0),
    .cp0_tlb_write_data_paddr_1(u_mips_cpu_cp0_tlb_write_data_paddr_1),
    .cp0_tlb_write_data_c_0(u_mips_cpu_cp0_tlb_write_data_c_0),
    .cp0_tlb_write_data_c_1(u_mips_cpu_cp0_tlb_write_data_c_1),
    .cp0_tlb_write_data_d_0(u_mips_cpu_cp0_tlb_write_data_d_0),
    .cp0_tlb_write_data_d_1(u_mips_cpu_cp0_tlb_write_data_d_1),
    .cp0_tlb_write_data_v_0(u_mips_cpu_cp0_tlb_write_data_v_0),
    .cp0_tlb_write_data_v_1(u_mips_cpu_cp0_tlb_write_data_v_1),
    .tlb_write_en(u_mips_cpu_tlb_write_en)
  );
  inst_cache inst_cache ( // @[my_cpu_top.scala 320:30]
    .clock(inst_cache_clock),
    .reset(inst_cache_reset),
    .io_port_araddr(inst_cache_io_port_araddr),
    .io_port_arlen(inst_cache_io_port_arlen),
    .io_port_arburst(inst_cache_io_port_arburst),
    .io_port_arvalid(inst_cache_io_port_arvalid),
    .io_port_arready(inst_cache_io_port_arready),
    .io_port_rdata(inst_cache_io_port_rdata),
    .io_port_rlast(inst_cache_io_port_rlast),
    .io_port_rvalid(inst_cache_io_port_rvalid),
    .io_port_sram_req(inst_cache_io_port_sram_req),
    .io_port_sram_addr(inst_cache_io_port_sram_addr),
    .io_port_sram_write_en(inst_cache_io_port_sram_write_en),
    .io_port_sram_rdata_L(inst_cache_io_port_sram_rdata_L),
    .io_port_sram_cache(inst_cache_io_port_sram_cache),
    .io_stage2_flush(inst_cache_io_stage2_flush),
    .io_stage2_stall(inst_cache_io_stage2_stall),
    .io_stage1_valid_flush(inst_cache_io_stage1_valid_flush),
    .io_inst_ready_to_use(inst_cache_io_inst_ready_to_use),
    .io_inst_buffer_full(inst_cache_io_inst_buffer_full),
    .io_stage2_exception(inst_cache_io_stage2_exception),
    .io_cp0_asid(inst_cache_io_cp0_asid),
    .io_v_addr_for_tlb(inst_cache_io_v_addr_for_tlb),
    .io_p_addr_for_tlb(inst_cache_io_p_addr_for_tlb),
    .io_tlb_req(inst_cache_io_tlb_req),
    .io_tlb_exception(inst_cache_io_tlb_exception),
    .io_inst_ready_branch(inst_cache_io_inst_ready_branch),
    .io_inst_buffer_empty(inst_cache_io_inst_buffer_empty)
  );
  data_cache data_cache ( // @[my_cpu_top.scala 322:30]
    .clock(data_cache_clock),
    .reset(data_cache_reset),
    .io_port_araddr(data_cache_io_port_araddr),
    .io_port_arlen(data_cache_io_port_arlen),
    .io_port_arsize(data_cache_io_port_arsize),
    .io_port_arburst(data_cache_io_port_arburst),
    .io_port_arvalid(data_cache_io_port_arvalid),
    .io_port_arready(data_cache_io_port_arready),
    .io_port_rdata(data_cache_io_port_rdata),
    .io_port_rlast(data_cache_io_port_rlast),
    .io_port_rvalid(data_cache_io_port_rvalid),
    .io_port_awaddr(data_cache_io_port_awaddr),
    .io_port_awlen(data_cache_io_port_awlen),
    .io_port_awsize(data_cache_io_port_awsize),
    .io_port_awburst(data_cache_io_port_awburst),
    .io_port_awvalid(data_cache_io_port_awvalid),
    .io_port_awready(data_cache_io_port_awready),
    .io_port_wdata(data_cache_io_port_wdata),
    .io_port_wstrb(data_cache_io_port_wstrb),
    .io_port_wlast(data_cache_io_port_wlast),
    .io_port_wvalid(data_cache_io_port_wvalid),
    .io_port_wready(data_cache_io_port_wready),
    .io_port_bvalid(data_cache_io_port_bvalid),
    .io_port_sram_req(data_cache_io_port_sram_req),
    .io_port_sram_wr(data_cache_io_port_sram_wr),
    .io_port_sram_size(data_cache_io_port_sram_size),
    .io_port_sram_addr(data_cache_io_port_sram_addr),
    .io_port_sram_wdata(data_cache_io_port_sram_wdata),
    .io_port_sram_rdata(data_cache_io_port_sram_rdata),
    .io_port_sram_cache(data_cache_io_port_sram_cache),
    .io_stage2_stall(data_cache_io_stage2_stall),
    .io_stage1_wr(data_cache_io_stage1_wr),
    .io_v_addr_for_tlb(data_cache_io_v_addr_for_tlb),
    .io_p_addr_for_tlb(data_cache_io_p_addr_for_tlb),
    .io_tlb_req(data_cache_io_tlb_req),
    .io_tlb_exception(data_cache_io_tlb_exception),
    .io_stage1_tlb_exception(data_cache_io_stage1_tlb_exception),
    .io_data_wstrb(data_cache_io_data_wstrb)
  );
  double_ports_tlb_for_inst_and_data double_ports_tlb_for_inst_and_data ( // @[my_cpu_top.scala 325:22]
    .clock(double_ports_tlb_for_inst_and_data_clock),
    .reset(double_ports_tlb_for_inst_and_data_reset),
    .io_cp0_asid(double_ports_tlb_for_inst_and_data_io_cp0_asid),
    .io_tlb_write_index(double_ports_tlb_for_inst_and_data_io_tlb_write_index),
    .io_tlb_read_index(double_ports_tlb_for_inst_and_data_io_tlb_read_index),
    .io_tlb_write_en(double_ports_tlb_for_inst_and_data_io_tlb_write_en),
    .io_tlb_search_index(double_ports_tlb_for_inst_and_data_io_tlb_search_index),
    .io_tlb_search_hit(double_ports_tlb_for_inst_and_data_io_tlb_search_hit),
    .io_tlb_dirty_exception(double_ports_tlb_for_inst_and_data_io_tlb_dirty_exception),
    .io_tlb_write_port_vaddr(double_ports_tlb_for_inst_and_data_io_tlb_write_port_vaddr),
    .io_tlb_write_port_asid(double_ports_tlb_for_inst_and_data_io_tlb_write_port_asid),
    .io_tlb_write_port_g(double_ports_tlb_for_inst_and_data_io_tlb_write_port_g),
    .io_tlb_write_port_paddr_0(double_ports_tlb_for_inst_and_data_io_tlb_write_port_paddr_0),
    .io_tlb_write_port_paddr_1(double_ports_tlb_for_inst_and_data_io_tlb_write_port_paddr_1),
    .io_tlb_write_port_c_0(double_ports_tlb_for_inst_and_data_io_tlb_write_port_c_0),
    .io_tlb_write_port_c_1(double_ports_tlb_for_inst_and_data_io_tlb_write_port_c_1),
    .io_tlb_write_port_d_0(double_ports_tlb_for_inst_and_data_io_tlb_write_port_d_0),
    .io_tlb_write_port_d_1(double_ports_tlb_for_inst_and_data_io_tlb_write_port_d_1),
    .io_tlb_write_port_v_0(double_ports_tlb_for_inst_and_data_io_tlb_write_port_v_0),
    .io_tlb_write_port_v_1(double_ports_tlb_for_inst_and_data_io_tlb_write_port_v_1),
    .io_tlb_read_port_vaddr(double_ports_tlb_for_inst_and_data_io_tlb_read_port_vaddr),
    .io_tlb_read_port_asid(double_ports_tlb_for_inst_and_data_io_tlb_read_port_asid),
    .io_tlb_read_port_g(double_ports_tlb_for_inst_and_data_io_tlb_read_port_g),
    .io_tlb_read_port_paddr_0(double_ports_tlb_for_inst_and_data_io_tlb_read_port_paddr_0),
    .io_tlb_read_port_paddr_1(double_ports_tlb_for_inst_and_data_io_tlb_read_port_paddr_1),
    .io_tlb_read_port_c_0(double_ports_tlb_for_inst_and_data_io_tlb_read_port_c_0),
    .io_tlb_read_port_c_1(double_ports_tlb_for_inst_and_data_io_tlb_read_port_c_1),
    .io_tlb_read_port_d_0(double_ports_tlb_for_inst_and_data_io_tlb_read_port_d_0),
    .io_tlb_read_port_d_1(double_ports_tlb_for_inst_and_data_io_tlb_read_port_d_1),
    .io_tlb_read_port_v_0(double_ports_tlb_for_inst_and_data_io_tlb_read_port_v_0),
    .io_tlb_read_port_v_1(double_ports_tlb_for_inst_and_data_io_tlb_read_port_v_1),
    .io_icache_port_vaddr(double_ports_tlb_for_inst_and_data_io_icache_port_vaddr),
    .io_icache_port_paddr(double_ports_tlb_for_inst_and_data_io_icache_port_paddr),
    .io_icache_port_req(double_ports_tlb_for_inst_and_data_io_icache_port_req),
    .io_icache_port_tlb_search_not_hit_exception(
      double_ports_tlb_for_inst_and_data_io_icache_port_tlb_search_not_hit_exception),
    .io_icache_port_tlb_search_ineffective_exception(
      double_ports_tlb_for_inst_and_data_io_icache_port_tlb_search_ineffective_exception),
    .io_dcache_port_vaddr(double_ports_tlb_for_inst_and_data_io_dcache_port_vaddr),
    .io_dcache_port_paddr(double_ports_tlb_for_inst_and_data_io_dcache_port_paddr),
    .io_dcache_port_req(double_ports_tlb_for_inst_and_data_io_dcache_port_req),
    .io_dcache_port_wr(double_ports_tlb_for_inst_and_data_io_dcache_port_wr),
    .io_dcache_port_tlb_search_not_hit_exception(
      double_ports_tlb_for_inst_and_data_io_dcache_port_tlb_search_not_hit_exception),
    .io_dcache_port_tlb_search_ineffective_exception(
      double_ports_tlb_for_inst_and_data_io_dcache_port_tlb_search_ineffective_exception)
  );
  assign arid = u_axi_cache_bridge_m_axi_arid; // @[my_cpu_top.scala 483:25]
  assign araddr = u_axi_cache_bridge_m_axi_araddr; // @[my_cpu_top.scala 484:25]
  assign arlen = u_axi_cache_bridge_m_axi_arlen; // @[my_cpu_top.scala 485:25]
  assign arsize = u_axi_cache_bridge_m_axi_arsize; // @[my_cpu_top.scala 486:25]
  assign arburst = u_axi_cache_bridge_m_axi_arburst; // @[my_cpu_top.scala 487:25]
  assign arlock = u_axi_cache_bridge_m_axi_arlock; // @[my_cpu_top.scala 488:25]
  assign arcache = u_axi_cache_bridge_m_axi_arcache; // @[my_cpu_top.scala 489:25]
  assign arprot = u_axi_cache_bridge_m_axi_arprot; // @[my_cpu_top.scala 490:25]
  assign arvalid = u_axi_cache_bridge_m_axi_arvalid; // @[my_cpu_top.scala 492:25]
  assign rready = u_axi_cache_bridge_m_axi_rready; // @[my_cpu_top.scala 500:25]
  assign awid = u_axi_cache_bridge_m_axi_awid; // @[my_cpu_top.scala 460:25]
  assign awaddr = u_axi_cache_bridge_m_axi_awaddr; // @[my_cpu_top.scala 461:25]
  assign awlen = u_axi_cache_bridge_m_axi_awlen; // @[my_cpu_top.scala 462:25]
  assign awsize = u_axi_cache_bridge_m_axi_awsize; // @[my_cpu_top.scala 463:25]
  assign awburst = u_axi_cache_bridge_m_axi_awburst; // @[my_cpu_top.scala 464:25]
  assign awlock = u_axi_cache_bridge_m_axi_awlock; // @[my_cpu_top.scala 465:25]
  assign awcache = u_axi_cache_bridge_m_axi_awcache; // @[my_cpu_top.scala 466:25]
  assign awprot = u_axi_cache_bridge_m_axi_awprot; // @[my_cpu_top.scala 467:25]
  assign awvalid = u_axi_cache_bridge_m_axi_awvalid; // @[my_cpu_top.scala 469:25]
  assign wid = u_axi_cache_bridge_m_axi_wid; // @[my_cpu_top.scala 472:45]
  assign wdata = u_axi_cache_bridge_m_axi_wdata; // @[my_cpu_top.scala 473:45]
  assign wstrb = u_axi_cache_bridge_m_axi_wstrb; // @[my_cpu_top.scala 474:45]
  assign wlast = u_axi_cache_bridge_m_axi_wlast; // @[my_cpu_top.scala 475:45]
  assign wvalid = u_axi_cache_bridge_m_axi_wvalid; // @[my_cpu_top.scala 476:45]
  assign bready = u_axi_cache_bridge_m_axi_bready; // @[my_cpu_top.scala 481:25]
  assign debug_wb_pc = u_mips_cpu_debug_wb_pc; // @[my_cpu_top.scala 384:29]
  assign debug_wb_rf_wen = u_mips_cpu_debug_wb_rf_wen; // @[my_cpu_top.scala 386:29]
  assign debug_wb_rf_wnum = u_mips_cpu_debug_wb_rf_wnum; // @[my_cpu_top.scala 387:29]
  assign debug_wb_rf_wdata = u_mips_cpu_debug_wb_rf_wdata; // @[my_cpu_top.scala 385:29]
  assign u_axi_cache_bridge_aclk = aclk; // @[my_cpu_top.scala 401:44]
  assign u_axi_cache_bridge_aresetn = aresetn; // @[my_cpu_top.scala 402:44]
  assign u_axi_cache_bridge_s_axi_awid = 8'h11; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_awaddr = {data_cache_io_port_awaddr,32'h0}; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_awlen = {data_cache_io_port_awlen,4'h0}; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_awsize = {data_cache_io_port_awsize,3'h2}; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_awburst = {data_cache_io_port_awburst,2'h0}; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_awlock = 4'h0; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_awcache = 8'h0; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_awprot = 6'h0; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_awqos = 8'h0; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_awvalid = {data_cache_io_port_awvalid,1'h0}; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_wid = 8'h11; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_wdata = {data_cache_io_port_wdata,32'h0}; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_wstrb = {data_cache_io_port_wstrb,4'h0}; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_wlast = {data_cache_io_port_wlast,1'h0}; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_wvalid = {data_cache_io_port_wvalid,1'h0}; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_bready = 2'h2; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_arid = 8'h10; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_araddr = {data_cache_io_port_araddr,inst_cache_io_port_araddr}; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_arlen = {data_cache_io_port_arlen,inst_cache_io_port_arlen}; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_arsize = {data_cache_io_port_arsize,3'h2}; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_arburst = {data_cache_io_port_arburst,inst_cache_io_port_arburst}; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_arlock = 4'h0; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_arcache = 8'h0; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_arprot = 6'h0; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_arqos = 8'h0; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_arvalid = {data_cache_io_port_arvalid,inst_cache_io_port_arvalid}; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_s_axi_rready = 2'h3; // @[Cat.scala 31:58]
  assign u_axi_cache_bridge_m_axi_awready = awready; // @[my_cpu_top.scala 471:45]
  assign u_axi_cache_bridge_m_axi_wready = wready; // @[my_cpu_top.scala 477:45]
  assign u_axi_cache_bridge_m_axi_bid = bid; // @[my_cpu_top.scala 478:45]
  assign u_axi_cache_bridge_m_axi_bresp = bresp; // @[my_cpu_top.scala 479:45]
  assign u_axi_cache_bridge_m_axi_bvalid = bvalid; // @[my_cpu_top.scala 480:45]
  assign u_axi_cache_bridge_m_axi_arready = arready; // @[my_cpu_top.scala 494:43]
  assign u_axi_cache_bridge_m_axi_rid = rid; // @[my_cpu_top.scala 495:40]
  assign u_axi_cache_bridge_m_axi_rdata = rdata; // @[my_cpu_top.scala 496:40]
  assign u_axi_cache_bridge_m_axi_rresp = rresp; // @[my_cpu_top.scala 497:40]
  assign u_axi_cache_bridge_m_axi_rlast = rlast; // @[my_cpu_top.scala 498:40]
  assign u_axi_cache_bridge_m_axi_rvalid = rvalid; // @[my_cpu_top.scala 499:40]
  assign u_mips_cpu_ext_int = ext_int; // @[my_cpu_top.scala 390:29]
  assign u_mips_cpu_resetn = aresetn; // @[my_cpu_top.scala 389:29]
  assign u_mips_cpu_clk = aclk; // @[my_cpu_top.scala 388:29]
  assign u_mips_cpu_inst_sram_rdata_L = inst_cache_io_port_sram_rdata_L; // @[my_cpu_top.scala 370:31]
  assign u_mips_cpu_inst_write_en = inst_cache_io_port_sram_write_en; // @[my_cpu_top.scala 378:30]
  assign u_mips_cpu_inst_tlb_exception = inst_cache_io_stage2_exception; // @[my_cpu_top.scala 380:35]
  assign u_mips_cpu_stage2_stall = inst_cache_io_stage2_stall; // @[my_cpu_top.scala 391:34]
  assign u_mips_cpu_data_sram_rdata = data_cache_io_port_sram_rdata; // @[my_cpu_top.scala 357:27]
  assign u_mips_cpu_data_stage2_stall = data_cache_io_stage2_stall; // @[my_cpu_top.scala 379:34]
  assign u_mips_cpu_data_tlb_exception = data_cache_io_stage1_tlb_exception; // @[my_cpu_top.scala 381:35]
  assign u_mips_cpu_tlb_search_index = double_ports_tlb_for_inst_and_data_io_tlb_search_index; // @[my_cpu_top.scala 394:33]
  assign u_mips_cpu_tlb_search_hit = double_ports_tlb_for_inst_and_data_io_tlb_search_hit; // @[my_cpu_top.scala 392:32]
  assign u_mips_cpu_cp0_tlb_write_data_vaddr = double_ports_tlb_for_inst_and_data_io_tlb_read_port_vaddr; // @[my_cpu_top.scala 395:35]
  assign u_mips_cpu_cp0_tlb_write_data_asid = double_ports_tlb_for_inst_and_data_io_tlb_read_port_asid; // @[my_cpu_top.scala 395:35]
  assign u_mips_cpu_cp0_tlb_write_data_g = double_ports_tlb_for_inst_and_data_io_tlb_read_port_g; // @[my_cpu_top.scala 395:35]
  assign u_mips_cpu_cp0_tlb_write_data_paddr_0 = double_ports_tlb_for_inst_and_data_io_tlb_read_port_paddr_0; // @[my_cpu_top.scala 395:35]
  assign u_mips_cpu_cp0_tlb_write_data_paddr_1 = double_ports_tlb_for_inst_and_data_io_tlb_read_port_paddr_1; // @[my_cpu_top.scala 395:35]
  assign u_mips_cpu_cp0_tlb_write_data_c_0 = double_ports_tlb_for_inst_and_data_io_tlb_read_port_c_0; // @[my_cpu_top.scala 395:35]
  assign u_mips_cpu_cp0_tlb_write_data_c_1 = double_ports_tlb_for_inst_and_data_io_tlb_read_port_c_1; // @[my_cpu_top.scala 395:35]
  assign u_mips_cpu_cp0_tlb_write_data_d_0 = double_ports_tlb_for_inst_and_data_io_tlb_read_port_d_0; // @[my_cpu_top.scala 395:35]
  assign u_mips_cpu_cp0_tlb_write_data_d_1 = double_ports_tlb_for_inst_and_data_io_tlb_read_port_d_1; // @[my_cpu_top.scala 395:35]
  assign u_mips_cpu_cp0_tlb_write_data_v_0 = double_ports_tlb_for_inst_and_data_io_tlb_read_port_v_0; // @[my_cpu_top.scala 395:35]
  assign u_mips_cpu_cp0_tlb_write_data_v_1 = double_ports_tlb_for_inst_and_data_io_tlb_read_port_v_1; // @[my_cpu_top.scala 395:35]
  assign inst_cache_clock = aclk; // @[my_cpu_top.scala 317:23]
  assign inst_cache_reset = ~aresetn; // @[my_cpu_top.scala 317:42]
  assign inst_cache_io_port_arready = u_axi_cache_bridge_s_axi_arready[0]; // @[my_cpu_top.scala 445:69]
  assign inst_cache_io_port_rdata = u_axi_cache_bridge_s_axi_rdata[31:0]; // @[my_cpu_top.scala 449:67]
  assign inst_cache_io_port_rlast = u_axi_cache_bridge_s_axi_rlast[0]; // @[my_cpu_top.scala 453:67]
  assign inst_cache_io_port_rvalid = u_axi_cache_bridge_s_axi_rvalid[0]; // @[my_cpu_top.scala 455:68]
  assign inst_cache_io_port_sram_req = u_mips_cpu_inst_sram_en; // @[my_cpu_top.scala 364:29]
  assign inst_cache_io_port_sram_addr = u_mips_cpu_inst_sram_addr; // @[my_cpu_top.scala 361:29]
  assign inst_cache_io_port_sram_cache = u_mips_cpu_inst_cache; // @[my_cpu_top.scala 363:29]
  assign inst_cache_io_stage2_flush = u_mips_cpu_stage2_flush; // @[my_cpu_top.scala 442:31]
  assign inst_cache_io_stage1_valid_flush = u_mips_cpu_stage1_valid_flush; // @[my_cpu_top.scala 502:37]
  assign inst_cache_io_inst_ready_to_use = u_mips_cpu_inst_ready_to_use; // @[my_cpu_top.scala 503:36]
  assign inst_cache_io_inst_buffer_full = u_mips_cpu_inst_buffer_full; // @[my_cpu_top.scala 504:37]
  assign inst_cache_io_cp0_asid = u_mips_cpu_cp0_asid; // @[my_cpu_top.scala 369:29]
  assign inst_cache_io_p_addr_for_tlb = double_ports_tlb_for_inst_and_data_io_icache_port_paddr; // @[my_cpu_top.scala 332:34]
  assign inst_cache_io_tlb_exception = {
    double_ports_tlb_for_inst_and_data_io_icache_port_tlb_search_ineffective_exception,
    double_ports_tlb_for_inst_and_data_io_icache_port_tlb_search_not_hit_exception}; // @[Cat.scala 31:58]
  assign inst_cache_io_inst_ready_branch = u_mips_cpu_inst_ready_branch; // @[my_cpu_top.scala 368:36]
  assign inst_cache_io_inst_buffer_empty = u_mips_cpu_inst_buffer_empty; // @[my_cpu_top.scala 367:36]
  assign data_cache_clock = aclk; // @[my_cpu_top.scala 317:23]
  assign data_cache_reset = ~aresetn; // @[my_cpu_top.scala 317:42]
  assign data_cache_io_port_arready = u_axi_cache_bridge_s_axi_arready[1]; // @[my_cpu_top.scala 444:69]
  assign data_cache_io_port_rdata = u_axi_cache_bridge_s_axi_rdata[63:32]; // @[my_cpu_top.scala 448:67]
  assign data_cache_io_port_rlast = u_axi_cache_bridge_s_axi_rlast[1]; // @[my_cpu_top.scala 452:67]
  assign data_cache_io_port_rvalid = u_axi_cache_bridge_s_axi_rvalid[1]; // @[my_cpu_top.scala 454:68]
  assign data_cache_io_port_awready = u_axi_cache_bridge_s_axi_awready[1]; // @[my_cpu_top.scala 413:83]
  assign data_cache_io_port_wready = u_axi_cache_bridge_s_axi_wready[1]; // @[my_cpu_top.scala 421:58]
  assign data_cache_io_port_bvalid = u_axi_cache_bridge_s_axi_bvalid[1]; // @[my_cpu_top.scala 427:58]
  assign data_cache_io_port_sram_req = u_mips_cpu_data_sram_en; // @[my_cpu_top.scala 353:23]
  assign data_cache_io_port_sram_wr = u_mips_cpu_data_sram_wen; // @[my_cpu_top.scala 354:23]
  assign data_cache_io_port_sram_size = u_mips_cpu_data_size; // @[my_cpu_top.scala 351:22]
  assign data_cache_io_port_sram_addr = u_mips_cpu_data_sram_addr; // @[my_cpu_top.scala 350:22]
  assign data_cache_io_port_sram_wdata = u_mips_cpu_data_sram_wdata; // @[my_cpu_top.scala 355:23]
  assign data_cache_io_port_sram_cache = u_mips_cpu_data_cache; // @[my_cpu_top.scala 352:23]
  assign data_cache_io_p_addr_for_tlb = double_ports_tlb_for_inst_and_data_io_dcache_port_paddr; // @[my_cpu_top.scala 341:33]
  assign data_cache_io_tlb_exception = {hi,
    double_ports_tlb_for_inst_and_data_io_dcache_port_tlb_search_not_hit_exception}; // @[Cat.scala 31:58]
  assign data_cache_io_data_wstrb = u_mips_cpu_data_wstrb; // @[my_cpu_top.scala 356:29]
  assign double_ports_tlb_for_inst_and_data_clock = aclk; // @[my_cpu_top.scala 317:23]
  assign double_ports_tlb_for_inst_and_data_reset = ~aresetn; // @[my_cpu_top.scala 317:42]
  assign double_ports_tlb_for_inst_and_data_io_cp0_asid = u_mips_cpu_cp0_asid; // @[my_cpu_top.scala 327:27]
  assign double_ports_tlb_for_inst_and_data_io_tlb_write_index = u_mips_cpu_tlb_write_index; // @[my_cpu_top.scala 398:26]
  assign double_ports_tlb_for_inst_and_data_io_tlb_read_index = u_mips_cpu_tlb_read_index; // @[my_cpu_top.scala 399:26]
  assign double_ports_tlb_for_inst_and_data_io_tlb_write_en = u_mips_cpu_tlb_write_en; // @[my_cpu_top.scala 396:26]
  assign double_ports_tlb_for_inst_and_data_io_tlb_write_port_vaddr = u_mips_cpu_cp0_tlb_read_data_vaddr; // @[my_cpu_top.scala 397:26]
  assign double_ports_tlb_for_inst_and_data_io_tlb_write_port_asid = u_mips_cpu_cp0_tlb_read_data_asid; // @[my_cpu_top.scala 397:26]
  assign double_ports_tlb_for_inst_and_data_io_tlb_write_port_g = u_mips_cpu_cp0_tlb_read_data_g; // @[my_cpu_top.scala 397:26]
  assign double_ports_tlb_for_inst_and_data_io_tlb_write_port_paddr_0 = u_mips_cpu_cp0_tlb_read_data_paddr_0; // @[my_cpu_top.scala 397:26]
  assign double_ports_tlb_for_inst_and_data_io_tlb_write_port_paddr_1 = u_mips_cpu_cp0_tlb_read_data_paddr_1; // @[my_cpu_top.scala 397:26]
  assign double_ports_tlb_for_inst_and_data_io_tlb_write_port_c_0 = u_mips_cpu_cp0_tlb_read_data_c_0; // @[my_cpu_top.scala 397:26]
  assign double_ports_tlb_for_inst_and_data_io_tlb_write_port_c_1 = u_mips_cpu_cp0_tlb_read_data_c_1; // @[my_cpu_top.scala 397:26]
  assign double_ports_tlb_for_inst_and_data_io_tlb_write_port_d_0 = u_mips_cpu_cp0_tlb_read_data_d_0; // @[my_cpu_top.scala 397:26]
  assign double_ports_tlb_for_inst_and_data_io_tlb_write_port_d_1 = u_mips_cpu_cp0_tlb_read_data_d_1; // @[my_cpu_top.scala 397:26]
  assign double_ports_tlb_for_inst_and_data_io_tlb_write_port_v_0 = u_mips_cpu_cp0_tlb_read_data_v_0; // @[my_cpu_top.scala 397:26]
  assign double_ports_tlb_for_inst_and_data_io_tlb_write_port_v_1 = u_mips_cpu_cp0_tlb_read_data_v_1; // @[my_cpu_top.scala 397:26]
  assign double_ports_tlb_for_inst_and_data_io_icache_port_vaddr = inst_cache_io_v_addr_for_tlb; // @[my_cpu_top.scala 328:27]
  assign double_ports_tlb_for_inst_and_data_io_icache_port_req = inst_cache_io_tlb_req; // @[my_cpu_top.scala 329:27]
  assign double_ports_tlb_for_inst_and_data_io_dcache_port_vaddr = u_mips_cpu_tlbp_search_en ?
    u_mips_cpu_tlbp_search_vaddr : data_cache_io_v_addr_for_tlb; // @[my_cpu_top.scala 338:33]
  assign double_ports_tlb_for_inst_and_data_io_dcache_port_req = data_cache_io_tlb_req; // @[my_cpu_top.scala 339:27]
  assign double_ports_tlb_for_inst_and_data_io_dcache_port_wr = data_cache_io_stage1_wr; // @[my_cpu_top.scala 340:27]
endmodule
